
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_ALU_ENTITY is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_ALU_ENTITY;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ALU_ENTITY.all;

entity ALU_ENTITY_DW02_mult_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  PRODUCT
         : out std_logic_vector (63 downto 0));

end ALU_ENTITY_DW02_mult_0;

architecture SYN_csa of ALU_ENTITY_DW02_mult_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal ab_31_0_port, ab_30_1_port, ab_30_0_port, ab_29_2_port, ab_29_1_port,
      ab_29_0_port, ab_28_3_port, ab_28_2_port, ab_28_1_port, ab_28_0_port, 
      ab_27_4_port, ab_27_3_port, ab_27_2_port, ab_27_1_port, ab_27_0_port, 
      ab_26_5_port, ab_26_4_port, ab_26_3_port, ab_26_2_port, ab_26_1_port, 
      ab_26_0_port, ab_25_6_port, ab_25_5_port, ab_25_4_port, ab_25_3_port, 
      ab_25_2_port, ab_25_1_port, ab_25_0_port, ab_24_7_port, ab_24_6_port, 
      ab_24_5_port, ab_24_4_port, ab_24_3_port, ab_24_2_port, ab_24_1_port, 
      ab_24_0_port, ab_23_8_port, ab_23_7_port, ab_23_6_port, ab_23_5_port, 
      ab_23_4_port, ab_23_3_port, ab_23_2_port, ab_23_1_port, ab_23_0_port, 
      ab_22_9_port, ab_22_8_port, ab_22_7_port, ab_22_6_port, ab_22_5_port, 
      ab_22_4_port, ab_22_3_port, ab_22_2_port, ab_22_1_port, ab_22_0_port, 
      ab_21_10_port, ab_21_9_port, ab_21_8_port, ab_21_7_port, ab_21_6_port, 
      ab_21_5_port, ab_21_4_port, ab_21_3_port, ab_21_2_port, ab_21_1_port, 
      ab_21_0_port, ab_20_11_port, ab_20_10_port, ab_20_9_port, ab_20_8_port, 
      ab_20_7_port, ab_20_6_port, ab_20_5_port, ab_20_4_port, ab_20_3_port, 
      ab_20_2_port, ab_20_1_port, ab_20_0_port, ab_19_12_port, ab_19_11_port, 
      ab_19_10_port, ab_19_9_port, ab_19_8_port, ab_19_7_port, ab_19_6_port, 
      ab_19_5_port, ab_19_4_port, ab_19_3_port, ab_19_2_port, ab_19_1_port, 
      ab_19_0_port, ab_18_13_port, ab_18_12_port, ab_18_11_port, ab_18_10_port,
      ab_18_9_port, ab_18_8_port, ab_18_7_port, ab_18_6_port, ab_18_5_port, 
      ab_18_4_port, ab_18_3_port, ab_18_2_port, ab_18_1_port, ab_18_0_port, 
      ab_17_14_port, ab_17_13_port, ab_17_12_port, ab_17_11_port, ab_17_10_port
      , ab_17_9_port, ab_17_8_port, ab_17_7_port, ab_17_6_port, ab_17_5_port, 
      ab_17_4_port, ab_17_3_port, ab_17_2_port, ab_17_1_port, ab_17_0_port, 
      ab_16_15_port, ab_16_14_port, ab_16_13_port, ab_16_12_port, ab_16_11_port
      , ab_16_10_port, ab_16_9_port, ab_16_8_port, ab_16_7_port, ab_16_6_port, 
      ab_16_5_port, ab_16_4_port, ab_16_3_port, ab_16_2_port, ab_16_1_port, 
      ab_16_0_port, ab_15_16_port, ab_15_15_port, ab_15_14_port, ab_15_13_port,
      ab_15_12_port, ab_15_11_port, ab_15_10_port, ab_15_9_port, ab_15_8_port, 
      ab_15_7_port, ab_15_6_port, ab_15_5_port, ab_15_4_port, ab_15_3_port, 
      ab_15_2_port, ab_15_1_port, ab_15_0_port, ab_14_17_port, ab_14_16_port, 
      ab_14_15_port, ab_14_14_port, ab_14_13_port, ab_14_12_port, ab_14_11_port
      , ab_14_10_port, ab_14_9_port, ab_14_8_port, ab_14_7_port, ab_14_6_port, 
      ab_14_5_port, ab_14_4_port, ab_14_3_port, ab_14_2_port, ab_14_1_port, 
      ab_14_0_port, ab_13_18_port, ab_13_17_port, ab_13_16_port, ab_13_15_port,
      ab_13_14_port, ab_13_13_port, ab_13_12_port, ab_13_11_port, ab_13_10_port
      , ab_13_9_port, ab_13_8_port, ab_13_7_port, ab_13_6_port, ab_13_5_port, 
      ab_13_4_port, ab_13_3_port, ab_13_2_port, ab_13_1_port, ab_13_0_port, 
      ab_12_19_port, ab_12_18_port, ab_12_17_port, ab_12_16_port, ab_12_15_port
      , ab_12_14_port, ab_12_13_port, ab_12_12_port, ab_12_11_port, 
      ab_12_10_port, ab_12_9_port, ab_12_8_port, ab_12_7_port, ab_12_6_port, 
      ab_12_5_port, ab_12_4_port, ab_12_3_port, ab_12_2_port, ab_12_1_port, 
      ab_12_0_port, ab_11_20_port, ab_11_19_port, ab_11_18_port, ab_11_17_port,
      ab_11_16_port, ab_11_15_port, ab_11_14_port, ab_11_13_port, ab_11_12_port
      , ab_11_11_port, ab_11_10_port, ab_11_9_port, ab_11_8_port, ab_11_7_port,
      ab_11_6_port, ab_11_5_port, ab_11_4_port, ab_11_3_port, ab_11_2_port, 
      ab_11_1_port, ab_11_0_port, ab_10_21_port, ab_10_20_port, ab_10_19_port, 
      ab_10_18_port, ab_10_17_port, ab_10_16_port, ab_10_15_port, ab_10_14_port
      , ab_10_13_port, ab_10_12_port, ab_10_11_port, ab_10_10_port, 
      ab_10_9_port, ab_10_8_port, ab_10_7_port, ab_10_6_port, ab_10_5_port, 
      ab_10_4_port, ab_10_3_port, ab_10_2_port, ab_10_1_port, ab_10_0_port, 
      ab_9_22_port, ab_9_21_port, ab_9_20_port, ab_9_19_port, ab_9_18_port, 
      ab_9_17_port, ab_9_16_port, ab_9_15_port, ab_9_14_port, ab_9_13_port, 
      ab_9_12_port, ab_9_11_port, ab_9_10_port, ab_9_9_port, ab_9_8_port, 
      ab_9_7_port, ab_9_6_port, ab_9_5_port, ab_9_4_port, ab_9_3_port, 
      ab_9_2_port, ab_9_1_port, ab_9_0_port, ab_8_23_port, ab_8_22_port, 
      ab_8_21_port, ab_8_20_port, ab_8_19_port, ab_8_18_port, ab_8_17_port, 
      ab_8_16_port, ab_8_15_port, ab_8_14_port, ab_8_13_port, ab_8_12_port, 
      ab_8_11_port, ab_8_10_port, ab_8_9_port, ab_8_8_port, ab_8_7_port, 
      ab_8_6_port, ab_8_5_port, ab_8_4_port, ab_8_3_port, ab_8_2_port, 
      ab_8_1_port, ab_8_0_port, ab_7_24_port, ab_7_23_port, ab_7_22_port, 
      ab_7_21_port, ab_7_20_port, ab_7_19_port, ab_7_18_port, ab_7_17_port, 
      ab_7_16_port, ab_7_15_port, ab_7_14_port, ab_7_13_port, ab_7_12_port, 
      ab_7_11_port, ab_7_10_port, ab_7_9_port, ab_7_8_port, ab_7_7_port, 
      ab_7_6_port, ab_7_5_port, ab_7_4_port, ab_7_3_port, ab_7_2_port, 
      ab_7_1_port, ab_7_0_port, ab_6_25_port, ab_6_24_port, ab_6_23_port, 
      ab_6_22_port, ab_6_21_port, ab_6_20_port, ab_6_19_port, ab_6_18_port, 
      ab_6_17_port, ab_6_16_port, ab_6_15_port, ab_6_14_port, ab_6_13_port, 
      ab_6_12_port, ab_6_11_port, ab_6_10_port, ab_6_9_port, ab_6_8_port, 
      ab_6_7_port, ab_6_6_port, ab_6_5_port, ab_6_4_port, ab_6_3_port, 
      ab_6_2_port, ab_6_1_port, ab_6_0_port, ab_5_26_port, ab_5_25_port, 
      ab_5_24_port, ab_5_23_port, ab_5_22_port, ab_5_21_port, ab_5_20_port, 
      ab_5_19_port, ab_5_18_port, ab_5_17_port, ab_5_16_port, ab_5_15_port, 
      ab_5_14_port, ab_5_13_port, ab_5_12_port, ab_5_11_port, ab_5_10_port, 
      ab_5_9_port, ab_5_8_port, ab_5_7_port, ab_5_6_port, ab_5_5_port, 
      ab_5_4_port, ab_5_3_port, ab_5_2_port, ab_5_1_port, ab_5_0_port, 
      ab_4_27_port, ab_4_26_port, ab_4_25_port, ab_4_24_port, ab_4_23_port, 
      ab_4_22_port, ab_4_21_port, ab_4_20_port, ab_4_19_port, ab_4_18_port, 
      ab_4_17_port, ab_4_16_port, ab_4_15_port, ab_4_14_port, ab_4_13_port, 
      ab_4_12_port, ab_4_11_port, ab_4_10_port, ab_4_9_port, ab_4_8_port, 
      ab_4_7_port, ab_4_6_port, ab_4_5_port, ab_4_4_port, ab_4_3_port, 
      ab_4_2_port, ab_4_1_port, ab_4_0_port, ab_3_28_port, ab_3_27_port, 
      ab_3_26_port, ab_3_25_port, ab_3_24_port, ab_3_23_port, ab_3_22_port, 
      ab_3_21_port, ab_3_20_port, ab_3_19_port, ab_3_18_port, ab_3_17_port, 
      ab_3_16_port, ab_3_15_port, ab_3_14_port, ab_3_13_port, ab_3_12_port, 
      ab_3_11_port, ab_3_10_port, ab_3_9_port, ab_3_8_port, ab_3_7_port, 
      ab_3_6_port, ab_3_5_port, ab_3_4_port, ab_3_3_port, ab_3_2_port, 
      ab_3_1_port, ab_3_0_port, ab_2_29_port, ab_2_28_port, ab_2_27_port, 
      ab_2_26_port, ab_2_25_port, ab_2_24_port, ab_2_23_port, ab_2_22_port, 
      ab_2_21_port, ab_2_20_port, ab_2_19_port, ab_2_18_port, ab_2_17_port, 
      ab_2_16_port, ab_2_15_port, ab_2_14_port, ab_2_13_port, ab_2_12_port, 
      ab_2_11_port, ab_2_10_port, ab_2_9_port, ab_2_8_port, ab_2_7_port, 
      ab_2_6_port, ab_2_5_port, ab_2_4_port, ab_2_3_port, ab_2_2_port, 
      ab_2_1_port, ab_2_0_port, ab_1_30_port, ab_1_29_port, ab_1_28_port, 
      ab_1_27_port, ab_1_26_port, ab_1_25_port, ab_1_24_port, ab_1_23_port, 
      ab_1_22_port, ab_1_21_port, ab_1_20_port, ab_1_19_port, ab_1_18_port, 
      ab_1_17_port, ab_1_16_port, ab_1_15_port, ab_1_14_port, ab_1_13_port, 
      ab_1_12_port, ab_1_11_port, ab_1_10_port, ab_1_9_port, ab_1_8_port, 
      ab_1_7_port, ab_1_6_port, ab_1_5_port, ab_1_4_port, ab_1_3_port, 
      ab_1_2_port, ab_1_1_port, ab_1_0_port, ab_0_31_port, ab_0_30_port, 
      ab_0_29_port, ab_0_28_port, ab_0_27_port, ab_0_26_port, ab_0_25_port, 
      ab_0_24_port, ab_0_23_port, ab_0_22_port, ab_0_21_port, ab_0_20_port, 
      ab_0_19_port, ab_0_18_port, ab_0_17_port, ab_0_16_port, ab_0_15_port, 
      ab_0_14_port, ab_0_13_port, ab_0_12_port, ab_0_11_port, ab_0_10_port, 
      ab_0_9_port, ab_0_8_port, ab_0_7_port, ab_0_6_port, ab_0_5_port, 
      ab_0_4_port, ab_0_3_port, ab_0_2_port, ab_0_1_port, CARRYB_15_15_port, 
      CARRYB_15_14_port, CARRYB_15_13_port, CARRYB_15_12_port, 
      CARRYB_15_11_port, CARRYB_15_10_port, CARRYB_15_9_port, CARRYB_15_8_port,
      CARRYB_15_7_port, CARRYB_15_6_port, CARRYB_15_5_port, CARRYB_15_4_port, 
      CARRYB_15_3_port, CARRYB_15_2_port, CARRYB_15_1_port, CARRYB_15_0_port, 
      CARRYB_14_16_port, CARRYB_14_15_port, CARRYB_14_14_port, 
      CARRYB_14_13_port, CARRYB_14_12_port, CARRYB_14_11_port, 
      CARRYB_14_10_port, CARRYB_14_9_port, CARRYB_14_8_port, CARRYB_14_7_port, 
      CARRYB_14_6_port, CARRYB_14_5_port, CARRYB_14_4_port, CARRYB_14_3_port, 
      CARRYB_14_2_port, CARRYB_14_1_port, CARRYB_14_0_port, CARRYB_13_17_port, 
      CARRYB_13_16_port, CARRYB_13_15_port, CARRYB_13_14_port, 
      CARRYB_13_13_port, CARRYB_13_12_port, CARRYB_13_11_port, 
      CARRYB_13_10_port, CARRYB_13_9_port, CARRYB_13_8_port, CARRYB_13_7_port, 
      CARRYB_13_6_port, CARRYB_13_5_port, CARRYB_13_4_port, CARRYB_13_3_port, 
      CARRYB_13_2_port, CARRYB_13_1_port, CARRYB_13_0_port, CARRYB_12_18_port, 
      CARRYB_12_17_port, CARRYB_12_16_port, CARRYB_12_15_port, 
      CARRYB_12_14_port, CARRYB_12_13_port, CARRYB_12_12_port, 
      CARRYB_12_11_port, CARRYB_12_10_port, CARRYB_12_9_port, CARRYB_12_8_port,
      CARRYB_12_7_port, CARRYB_12_6_port, CARRYB_12_5_port, CARRYB_12_4_port, 
      CARRYB_12_3_port, CARRYB_12_2_port, CARRYB_12_1_port, CARRYB_12_0_port, 
      CARRYB_11_19_port, CARRYB_11_18_port, CARRYB_11_17_port, 
      CARRYB_11_16_port, CARRYB_11_15_port, CARRYB_11_14_port, 
      CARRYB_11_13_port, CARRYB_11_12_port, CARRYB_11_11_port, 
      CARRYB_11_10_port, CARRYB_11_9_port, CARRYB_11_8_port, CARRYB_11_7_port, 
      CARRYB_11_6_port, CARRYB_11_5_port, CARRYB_11_4_port, CARRYB_11_3_port, 
      CARRYB_11_2_port, CARRYB_11_1_port, CARRYB_11_0_port, CARRYB_10_20_port, 
      CARRYB_10_19_port, CARRYB_10_18_port, CARRYB_10_17_port, 
      CARRYB_10_16_port, CARRYB_10_15_port, CARRYB_10_14_port, 
      CARRYB_10_13_port, CARRYB_10_12_port, CARRYB_10_11_port, 
      CARRYB_10_10_port, CARRYB_10_9_port, CARRYB_10_8_port, CARRYB_10_7_port, 
      CARRYB_10_6_port, CARRYB_10_5_port, CARRYB_10_4_port, CARRYB_10_3_port, 
      CARRYB_10_2_port, CARRYB_10_1_port, CARRYB_10_0_port, CARRYB_9_21_port, 
      CARRYB_9_20_port, CARRYB_9_19_port, CARRYB_9_18_port, CARRYB_9_17_port, 
      CARRYB_9_16_port, CARRYB_9_15_port, CARRYB_9_14_port, CARRYB_9_13_port, 
      CARRYB_9_12_port, CARRYB_9_11_port, CARRYB_9_10_port, CARRYB_9_9_port, 
      CARRYB_9_8_port, CARRYB_9_7_port, CARRYB_9_6_port, CARRYB_9_5_port, 
      CARRYB_9_4_port, CARRYB_9_3_port, CARRYB_9_2_port, CARRYB_9_1_port, 
      CARRYB_9_0_port, CARRYB_8_22_port, CARRYB_8_21_port, CARRYB_8_20_port, 
      CARRYB_8_19_port, CARRYB_8_18_port, CARRYB_8_17_port, CARRYB_8_16_port, 
      CARRYB_8_15_port, CARRYB_8_14_port, CARRYB_8_13_port, CARRYB_8_12_port, 
      CARRYB_8_11_port, CARRYB_8_10_port, CARRYB_8_9_port, CARRYB_8_8_port, 
      CARRYB_8_7_port, CARRYB_8_6_port, CARRYB_8_5_port, CARRYB_8_4_port, 
      CARRYB_8_3_port, CARRYB_8_2_port, CARRYB_8_1_port, CARRYB_8_0_port, 
      CARRYB_7_23_port, CARRYB_7_22_port, CARRYB_7_21_port, CARRYB_7_20_port, 
      CARRYB_7_19_port, CARRYB_7_18_port, CARRYB_7_17_port, CARRYB_7_16_port, 
      CARRYB_7_15_port, CARRYB_7_14_port, CARRYB_7_13_port, CARRYB_7_12_port, 
      CARRYB_7_11_port, CARRYB_7_10_port, CARRYB_7_9_port, CARRYB_7_8_port, 
      CARRYB_7_7_port, CARRYB_7_6_port, CARRYB_7_5_port, CARRYB_7_4_port, 
      CARRYB_7_3_port, CARRYB_7_2_port, CARRYB_7_1_port, CARRYB_7_0_port, 
      CARRYB_6_24_port, CARRYB_6_23_port, CARRYB_6_22_port, CARRYB_6_21_port, 
      CARRYB_6_20_port, CARRYB_6_19_port, CARRYB_6_18_port, CARRYB_6_17_port, 
      CARRYB_6_16_port, CARRYB_6_15_port, CARRYB_6_14_port, CARRYB_6_13_port, 
      CARRYB_6_12_port, CARRYB_6_11_port, CARRYB_6_10_port, CARRYB_6_9_port, 
      CARRYB_6_8_port, CARRYB_6_7_port, CARRYB_6_6_port, CARRYB_6_5_port, 
      CARRYB_6_4_port, CARRYB_6_3_port, CARRYB_6_2_port, CARRYB_6_1_port, 
      CARRYB_6_0_port, CARRYB_5_25_port, CARRYB_5_24_port, CARRYB_5_23_port, 
      CARRYB_5_22_port, CARRYB_5_21_port, CARRYB_5_20_port, CARRYB_5_19_port, 
      CARRYB_5_18_port, CARRYB_5_17_port, CARRYB_5_16_port, CARRYB_5_15_port, 
      CARRYB_5_14_port, CARRYB_5_13_port, CARRYB_5_12_port, CARRYB_5_11_port, 
      CARRYB_5_10_port, CARRYB_5_9_port, CARRYB_5_8_port, CARRYB_5_7_port, 
      CARRYB_5_6_port, CARRYB_5_5_port, CARRYB_5_4_port, CARRYB_5_3_port, 
      CARRYB_5_2_port, CARRYB_5_1_port, CARRYB_5_0_port, CARRYB_4_26_port, 
      CARRYB_4_25_port, CARRYB_4_24_port, CARRYB_4_23_port, CARRYB_4_22_port, 
      CARRYB_4_21_port, CARRYB_4_20_port, CARRYB_4_19_port, CARRYB_4_18_port, 
      CARRYB_4_17_port, CARRYB_4_16_port, CARRYB_4_15_port, CARRYB_4_14_port, 
      CARRYB_4_13_port, CARRYB_4_12_port, CARRYB_4_11_port, CARRYB_4_10_port, 
      CARRYB_4_9_port, CARRYB_4_8_port, CARRYB_4_7_port, CARRYB_4_6_port, 
      CARRYB_4_5_port, CARRYB_4_4_port, CARRYB_4_3_port, CARRYB_4_2_port, 
      CARRYB_4_1_port, CARRYB_4_0_port, CARRYB_3_27_port, CARRYB_3_26_port, 
      CARRYB_3_25_port, CARRYB_3_24_port, CARRYB_3_23_port, CARRYB_3_22_port, 
      CARRYB_3_21_port, CARRYB_3_20_port, CARRYB_3_19_port, CARRYB_3_18_port, 
      CARRYB_3_17_port, CARRYB_3_16_port, CARRYB_3_15_port, CARRYB_3_14_port, 
      CARRYB_3_13_port, CARRYB_3_12_port, CARRYB_3_11_port, CARRYB_3_10_port, 
      CARRYB_3_9_port, CARRYB_3_8_port, CARRYB_3_7_port, CARRYB_3_6_port, 
      CARRYB_3_5_port, CARRYB_3_4_port, CARRYB_3_3_port, CARRYB_3_2_port, 
      CARRYB_3_1_port, CARRYB_3_0_port, CARRYB_2_28_port, CARRYB_2_27_port, 
      CARRYB_2_26_port, CARRYB_2_25_port, CARRYB_2_24_port, CARRYB_2_23_port, 
      CARRYB_2_22_port, CARRYB_2_21_port, CARRYB_2_20_port, CARRYB_2_19_port, 
      CARRYB_2_18_port, CARRYB_2_17_port, CARRYB_2_16_port, CARRYB_2_15_port, 
      CARRYB_2_14_port, CARRYB_2_13_port, CARRYB_2_12_port, CARRYB_2_11_port, 
      CARRYB_2_10_port, CARRYB_2_9_port, CARRYB_2_8_port, CARRYB_2_7_port, 
      CARRYB_2_6_port, CARRYB_2_5_port, CARRYB_2_4_port, CARRYB_2_3_port, 
      CARRYB_2_2_port, CARRYB_2_1_port, CARRYB_2_0_port, SUMB_15_16_port, 
      SUMB_15_15_port, SUMB_15_14_port, SUMB_15_13_port, SUMB_15_12_port, 
      SUMB_15_11_port, SUMB_15_10_port, SUMB_15_9_port, SUMB_15_8_port, 
      SUMB_15_7_port, SUMB_15_6_port, SUMB_15_5_port, SUMB_15_4_port, 
      SUMB_15_3_port, SUMB_15_2_port, SUMB_15_1_port, SUMB_14_17_port, 
      SUMB_14_16_port, SUMB_14_15_port, SUMB_14_14_port, SUMB_14_13_port, 
      SUMB_14_12_port, SUMB_14_11_port, SUMB_14_10_port, SUMB_14_9_port, 
      SUMB_14_8_port, SUMB_14_7_port, SUMB_14_6_port, SUMB_14_5_port, 
      SUMB_14_4_port, SUMB_14_3_port, SUMB_14_2_port, SUMB_14_1_port, 
      SUMB_13_18_port, SUMB_13_17_port, SUMB_13_16_port, SUMB_13_15_port, 
      SUMB_13_14_port, SUMB_13_13_port, SUMB_13_12_port, SUMB_13_11_port, 
      SUMB_13_10_port, SUMB_13_9_port, SUMB_13_8_port, SUMB_13_7_port, 
      SUMB_13_6_port, SUMB_13_5_port, SUMB_13_4_port, SUMB_13_3_port, 
      SUMB_13_2_port, SUMB_13_1_port, SUMB_12_19_port, SUMB_12_18_port, 
      SUMB_12_17_port, SUMB_12_16_port, SUMB_12_15_port, SUMB_12_14_port, 
      SUMB_12_13_port, SUMB_12_12_port, SUMB_12_11_port, SUMB_12_10_port, 
      SUMB_12_9_port, SUMB_12_8_port, SUMB_12_7_port, SUMB_12_6_port, 
      SUMB_12_5_port, SUMB_12_4_port, SUMB_12_3_port, SUMB_12_2_port, 
      SUMB_12_1_port, SUMB_11_20_port, SUMB_11_19_port, SUMB_11_18_port, 
      SUMB_11_17_port, SUMB_11_16_port, SUMB_11_15_port, SUMB_11_14_port, 
      SUMB_11_13_port, SUMB_11_12_port, SUMB_11_11_port, SUMB_11_10_port, 
      SUMB_11_9_port, SUMB_11_8_port, SUMB_11_7_port, SUMB_11_6_port, 
      SUMB_11_5_port, SUMB_11_4_port, SUMB_11_3_port, SUMB_11_2_port, 
      SUMB_11_1_port, SUMB_10_21_port, SUMB_10_20_port, SUMB_10_19_port, 
      SUMB_10_18_port, SUMB_10_17_port, SUMB_10_16_port, SUMB_10_15_port, 
      SUMB_10_14_port, SUMB_10_13_port, SUMB_10_12_port, SUMB_10_11_port, 
      SUMB_10_10_port, SUMB_10_9_port, SUMB_10_8_port, SUMB_10_7_port, 
      SUMB_10_6_port, SUMB_10_5_port, SUMB_10_4_port, SUMB_10_3_port, 
      SUMB_10_2_port, SUMB_10_1_port, SUMB_9_22_port, SUMB_9_21_port, 
      SUMB_9_20_port, SUMB_9_19_port, SUMB_9_18_port, SUMB_9_17_port, 
      SUMB_9_16_port, SUMB_9_15_port, SUMB_9_14_port, SUMB_9_13_port, 
      SUMB_9_12_port, SUMB_9_11_port, SUMB_9_10_port, SUMB_9_9_port, 
      SUMB_9_8_port, SUMB_9_7_port, SUMB_9_6_port, SUMB_9_5_port, SUMB_9_4_port
      , SUMB_9_3_port, SUMB_9_2_port, SUMB_9_1_port, SUMB_8_23_port, 
      SUMB_8_22_port, SUMB_8_21_port, SUMB_8_20_port, SUMB_8_19_port, 
      SUMB_8_18_port, SUMB_8_17_port, SUMB_8_16_port, SUMB_8_15_port, 
      SUMB_8_14_port, SUMB_8_13_port, SUMB_8_12_port, SUMB_8_11_port, 
      SUMB_8_10_port, SUMB_8_9_port, SUMB_8_8_port, SUMB_8_7_port, 
      SUMB_8_6_port, SUMB_8_5_port, SUMB_8_4_port, SUMB_8_3_port, SUMB_8_2_port
      , SUMB_8_1_port, SUMB_7_24_port, SUMB_7_23_port, SUMB_7_22_port, 
      SUMB_7_21_port, SUMB_7_20_port, SUMB_7_19_port, SUMB_7_18_port, 
      SUMB_7_17_port, SUMB_7_16_port, SUMB_7_15_port, SUMB_7_14_port, 
      SUMB_7_13_port, SUMB_7_12_port, SUMB_7_11_port, SUMB_7_10_port, 
      SUMB_7_9_port, SUMB_7_8_port, SUMB_7_7_port, SUMB_7_6_port, SUMB_7_5_port
      , SUMB_7_4_port, SUMB_7_3_port, SUMB_7_2_port, SUMB_7_1_port, 
      SUMB_6_25_port, SUMB_6_24_port, SUMB_6_23_port, SUMB_6_22_port, 
      SUMB_6_21_port, SUMB_6_20_port, SUMB_6_19_port, SUMB_6_18_port, 
      SUMB_6_17_port, SUMB_6_16_port, SUMB_6_15_port, SUMB_6_14_port, 
      SUMB_6_13_port, SUMB_6_12_port, SUMB_6_11_port, SUMB_6_10_port, 
      SUMB_6_9_port, SUMB_6_8_port, SUMB_6_7_port, SUMB_6_6_port, SUMB_6_5_port
      , SUMB_6_4_port, SUMB_6_3_port, SUMB_6_2_port, SUMB_6_1_port, 
      SUMB_5_26_port, SUMB_5_25_port, SUMB_5_24_port, SUMB_5_23_port, 
      SUMB_5_22_port, SUMB_5_21_port, SUMB_5_20_port, SUMB_5_19_port, 
      SUMB_5_18_port, SUMB_5_17_port, SUMB_5_16_port, SUMB_5_15_port, 
      SUMB_5_14_port, SUMB_5_13_port, SUMB_5_12_port, SUMB_5_11_port, 
      SUMB_5_10_port, SUMB_5_9_port, SUMB_5_8_port, SUMB_5_7_port, 
      SUMB_5_6_port, SUMB_5_5_port, SUMB_5_4_port, SUMB_5_3_port, SUMB_5_2_port
      , SUMB_5_1_port, SUMB_4_27_port, SUMB_4_26_port, SUMB_4_25_port, 
      SUMB_4_24_port, SUMB_4_23_port, SUMB_4_22_port, SUMB_4_21_port, 
      SUMB_4_20_port, SUMB_4_19_port, SUMB_4_18_port, SUMB_4_17_port, 
      SUMB_4_16_port, SUMB_4_15_port, SUMB_4_14_port, SUMB_4_13_port, 
      SUMB_4_12_port, SUMB_4_11_port, SUMB_4_10_port, SUMB_4_9_port, 
      SUMB_4_8_port, SUMB_4_7_port, SUMB_4_6_port, SUMB_4_5_port, SUMB_4_4_port
      , SUMB_4_3_port, SUMB_4_2_port, SUMB_4_1_port, SUMB_3_28_port, 
      SUMB_3_27_port, SUMB_3_26_port, SUMB_3_25_port, SUMB_3_24_port, 
      SUMB_3_23_port, SUMB_3_22_port, SUMB_3_21_port, SUMB_3_20_port, 
      SUMB_3_19_port, SUMB_3_18_port, SUMB_3_17_port, SUMB_3_16_port, 
      SUMB_3_15_port, SUMB_3_14_port, SUMB_3_13_port, SUMB_3_12_port, 
      SUMB_3_11_port, SUMB_3_10_port, SUMB_3_9_port, SUMB_3_8_port, 
      SUMB_3_7_port, SUMB_3_6_port, SUMB_3_5_port, SUMB_3_4_port, SUMB_3_3_port
      , SUMB_3_2_port, SUMB_3_1_port, SUMB_2_29_port, SUMB_2_28_port, 
      SUMB_2_27_port, SUMB_2_26_port, SUMB_2_25_port, SUMB_2_24_port, 
      SUMB_2_23_port, SUMB_2_22_port, SUMB_2_21_port, SUMB_2_20_port, 
      SUMB_2_19_port, SUMB_2_18_port, SUMB_2_17_port, SUMB_2_16_port, 
      SUMB_2_15_port, SUMB_2_14_port, SUMB_2_13_port, SUMB_2_12_port, 
      SUMB_2_11_port, SUMB_2_10_port, SUMB_2_9_port, SUMB_2_8_port, 
      SUMB_2_7_port, SUMB_2_6_port, SUMB_2_5_port, SUMB_2_4_port, SUMB_2_3_port
      , SUMB_2_2_port, SUMB_2_1_port, CARRYB_30_0_port, CARRYB_29_1_port, 
      CARRYB_29_0_port, CARRYB_28_2_port, CARRYB_28_1_port, CARRYB_28_0_port, 
      CARRYB_27_3_port, CARRYB_27_2_port, CARRYB_27_1_port, CARRYB_27_0_port, 
      CARRYB_26_4_port, CARRYB_26_3_port, CARRYB_26_2_port, CARRYB_26_1_port, 
      CARRYB_26_0_port, CARRYB_25_5_port, CARRYB_25_4_port, CARRYB_25_3_port, 
      CARRYB_25_2_port, CARRYB_25_1_port, CARRYB_25_0_port, CARRYB_24_6_port, 
      CARRYB_24_5_port, CARRYB_24_4_port, CARRYB_24_3_port, CARRYB_24_2_port, 
      CARRYB_24_1_port, CARRYB_24_0_port, CARRYB_23_7_port, CARRYB_23_6_port, 
      CARRYB_23_5_port, CARRYB_23_4_port, CARRYB_23_3_port, CARRYB_23_2_port, 
      CARRYB_23_1_port, CARRYB_23_0_port, CARRYB_22_8_port, CARRYB_22_7_port, 
      CARRYB_22_6_port, CARRYB_22_5_port, CARRYB_22_4_port, CARRYB_22_3_port, 
      CARRYB_22_2_port, CARRYB_22_1_port, CARRYB_22_0_port, CARRYB_21_9_port, 
      CARRYB_21_8_port, CARRYB_21_7_port, CARRYB_21_6_port, CARRYB_21_5_port, 
      CARRYB_21_4_port, CARRYB_21_3_port, CARRYB_21_2_port, CARRYB_21_1_port, 
      CARRYB_21_0_port, CARRYB_20_10_port, CARRYB_20_9_port, CARRYB_20_8_port, 
      CARRYB_20_7_port, CARRYB_20_6_port, CARRYB_20_5_port, CARRYB_20_4_port, 
      CARRYB_20_3_port, CARRYB_20_2_port, CARRYB_20_1_port, CARRYB_20_0_port, 
      CARRYB_19_11_port, CARRYB_19_10_port, CARRYB_19_9_port, CARRYB_19_8_port,
      CARRYB_19_7_port, CARRYB_19_6_port, CARRYB_19_5_port, CARRYB_19_4_port, 
      CARRYB_19_3_port, CARRYB_19_2_port, CARRYB_19_1_port, CARRYB_19_0_port, 
      CARRYB_18_12_port, CARRYB_18_11_port, CARRYB_18_10_port, CARRYB_18_9_port
      , CARRYB_18_8_port, CARRYB_18_7_port, CARRYB_18_6_port, CARRYB_18_5_port,
      CARRYB_18_4_port, CARRYB_18_3_port, CARRYB_18_2_port, CARRYB_18_1_port, 
      CARRYB_18_0_port, CARRYB_17_13_port, CARRYB_17_12_port, CARRYB_17_11_port
      , CARRYB_17_10_port, CARRYB_17_9_port, CARRYB_17_8_port, CARRYB_17_7_port
      , CARRYB_17_6_port, CARRYB_17_5_port, CARRYB_17_4_port, CARRYB_17_3_port,
      CARRYB_17_2_port, CARRYB_17_1_port, CARRYB_17_0_port, CARRYB_16_14_port, 
      CARRYB_16_13_port, CARRYB_16_12_port, CARRYB_16_11_port, 
      CARRYB_16_10_port, CARRYB_16_9_port, CARRYB_16_8_port, CARRYB_16_7_port, 
      CARRYB_16_6_port, CARRYB_16_5_port, CARRYB_16_4_port, CARRYB_16_3_port, 
      CARRYB_16_2_port, CARRYB_16_1_port, CARRYB_16_0_port, SUMB_30_1_port, 
      SUMB_29_2_port, SUMB_29_1_port, SUMB_28_3_port, SUMB_28_2_port, 
      SUMB_28_1_port, SUMB_27_4_port, SUMB_27_3_port, SUMB_27_2_port, 
      SUMB_27_1_port, SUMB_26_5_port, SUMB_26_4_port, SUMB_26_3_port, 
      SUMB_26_2_port, SUMB_26_1_port, SUMB_25_6_port, SUMB_25_5_port, 
      SUMB_25_4_port, SUMB_25_3_port, SUMB_25_2_port, SUMB_25_1_port, 
      SUMB_24_7_port, SUMB_24_6_port, SUMB_24_5_port, SUMB_24_4_port, 
      SUMB_24_3_port, SUMB_24_2_port, SUMB_24_1_port, SUMB_23_8_port, 
      SUMB_23_7_port, SUMB_23_6_port, SUMB_23_5_port, SUMB_23_4_port, 
      SUMB_23_3_port, SUMB_23_2_port, SUMB_23_1_port, SUMB_22_9_port, 
      SUMB_22_8_port, SUMB_22_7_port, SUMB_22_6_port, SUMB_22_5_port, 
      SUMB_22_4_port, SUMB_22_3_port, SUMB_22_2_port, SUMB_22_1_port, 
      SUMB_21_10_port, SUMB_21_9_port, SUMB_21_8_port, SUMB_21_7_port, 
      SUMB_21_6_port, SUMB_21_5_port, SUMB_21_4_port, SUMB_21_3_port, 
      SUMB_21_2_port, SUMB_21_1_port, SUMB_20_11_port, SUMB_20_10_port, 
      SUMB_20_9_port, SUMB_20_8_port, SUMB_20_7_port, SUMB_20_6_port, 
      SUMB_20_5_port, SUMB_20_4_port, SUMB_20_3_port, SUMB_20_2_port, 
      SUMB_20_1_port, SUMB_19_12_port, SUMB_19_11_port, SUMB_19_10_port, 
      SUMB_19_9_port, SUMB_19_8_port, SUMB_19_7_port, SUMB_19_6_port, 
      SUMB_19_5_port, SUMB_19_4_port, SUMB_19_3_port, SUMB_19_2_port, 
      SUMB_19_1_port, SUMB_18_13_port, SUMB_18_12_port, SUMB_18_11_port, 
      SUMB_18_10_port, SUMB_18_9_port, SUMB_18_8_port, SUMB_18_7_port, 
      SUMB_18_6_port, SUMB_18_5_port, SUMB_18_4_port, SUMB_18_3_port, 
      SUMB_18_2_port, SUMB_18_1_port, SUMB_17_14_port, SUMB_17_13_port, 
      SUMB_17_12_port, SUMB_17_11_port, SUMB_17_10_port, SUMB_17_9_port, 
      SUMB_17_8_port, SUMB_17_7_port, SUMB_17_6_port, SUMB_17_5_port, 
      SUMB_17_4_port, SUMB_17_3_port, SUMB_17_2_port, SUMB_17_1_port, 
      SUMB_16_15_port, SUMB_16_14_port, SUMB_16_13_port, SUMB_16_12_port, 
      SUMB_16_11_port, SUMB_16_10_port, SUMB_16_9_port, SUMB_16_8_port, 
      SUMB_16_7_port, SUMB_16_6_port, SUMB_16_5_port, SUMB_16_4_port, 
      SUMB_16_3_port, SUMB_16_2_port, SUMB_16_1_port, n2, n3, n4, n5, n6, n7, 
      n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, 
      n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37
      , n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, 
      n52, n53, n54, n55, n56, n57, n58, n59, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n_1033, n_1034, n_1035, 
      n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, 
      n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, 
      n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062 : 
      std_logic;

begin
   
   S4_0 : FA_X1 port map( A => ab_31_0_port, B => CARRYB_30_0_port, CI => 
                           SUMB_30_1_port, CO => n_1033, S => PRODUCT(31));
   S1_30_0 : FA_X1 port map( A => ab_30_0_port, B => CARRYB_29_0_port, CI => 
                           SUMB_29_1_port, CO => CARRYB_30_0_port, S => 
                           PRODUCT(30));
   S2_30_1 : FA_X1 port map( A => ab_30_1_port, B => CARRYB_29_1_port, CI => 
                           SUMB_29_2_port, CO => n_1034, S => SUMB_30_1_port);
   S1_29_0 : FA_X1 port map( A => ab_29_0_port, B => CARRYB_28_0_port, CI => 
                           SUMB_28_1_port, CO => CARRYB_29_0_port, S => 
                           PRODUCT(29));
   S2_29_1 : FA_X1 port map( A => ab_29_1_port, B => CARRYB_28_1_port, CI => 
                           SUMB_28_2_port, CO => CARRYB_29_1_port, S => 
                           SUMB_29_1_port);
   S2_29_2 : FA_X1 port map( A => ab_29_2_port, B => CARRYB_28_2_port, CI => 
                           SUMB_28_3_port, CO => n_1035, S => SUMB_29_2_port);
   S1_28_0 : FA_X1 port map( A => ab_28_0_port, B => CARRYB_27_0_port, CI => 
                           SUMB_27_1_port, CO => CARRYB_28_0_port, S => 
                           PRODUCT(28));
   S2_28_1 : FA_X1 port map( A => ab_28_1_port, B => CARRYB_27_1_port, CI => 
                           SUMB_27_2_port, CO => CARRYB_28_1_port, S => 
                           SUMB_28_1_port);
   S2_28_2 : FA_X1 port map( A => ab_28_2_port, B => CARRYB_27_2_port, CI => 
                           SUMB_27_3_port, CO => CARRYB_28_2_port, S => 
                           SUMB_28_2_port);
   S2_28_3 : FA_X1 port map( A => ab_28_3_port, B => CARRYB_27_3_port, CI => 
                           SUMB_27_4_port, CO => n_1036, S => SUMB_28_3_port);
   S1_27_0 : FA_X1 port map( A => ab_27_0_port, B => CARRYB_26_0_port, CI => 
                           SUMB_26_1_port, CO => CARRYB_27_0_port, S => 
                           PRODUCT(27));
   S2_27_1 : FA_X1 port map( A => ab_27_1_port, B => CARRYB_26_1_port, CI => 
                           SUMB_26_2_port, CO => CARRYB_27_1_port, S => 
                           SUMB_27_1_port);
   S2_27_2 : FA_X1 port map( A => ab_27_2_port, B => CARRYB_26_2_port, CI => 
                           SUMB_26_3_port, CO => CARRYB_27_2_port, S => 
                           SUMB_27_2_port);
   S2_27_3 : FA_X1 port map( A => ab_27_3_port, B => CARRYB_26_3_port, CI => 
                           SUMB_26_4_port, CO => CARRYB_27_3_port, S => 
                           SUMB_27_3_port);
   S2_27_4 : FA_X1 port map( A => ab_27_4_port, B => CARRYB_26_4_port, CI => 
                           SUMB_26_5_port, CO => n_1037, S => SUMB_27_4_port);
   S1_26_0 : FA_X1 port map( A => ab_26_0_port, B => CARRYB_25_0_port, CI => 
                           SUMB_25_1_port, CO => CARRYB_26_0_port, S => 
                           PRODUCT(26));
   S2_26_1 : FA_X1 port map( A => ab_26_1_port, B => CARRYB_25_1_port, CI => 
                           SUMB_25_2_port, CO => CARRYB_26_1_port, S => 
                           SUMB_26_1_port);
   S2_26_2 : FA_X1 port map( A => ab_26_2_port, B => CARRYB_25_2_port, CI => 
                           SUMB_25_3_port, CO => CARRYB_26_2_port, S => 
                           SUMB_26_2_port);
   S2_26_3 : FA_X1 port map( A => ab_26_3_port, B => CARRYB_25_3_port, CI => 
                           SUMB_25_4_port, CO => CARRYB_26_3_port, S => 
                           SUMB_26_3_port);
   S2_26_4 : FA_X1 port map( A => ab_26_4_port, B => CARRYB_25_4_port, CI => 
                           SUMB_25_5_port, CO => CARRYB_26_4_port, S => 
                           SUMB_26_4_port);
   S2_26_5 : FA_X1 port map( A => ab_26_5_port, B => CARRYB_25_5_port, CI => 
                           SUMB_25_6_port, CO => n_1038, S => SUMB_26_5_port);
   S1_25_0 : FA_X1 port map( A => ab_25_0_port, B => CARRYB_24_0_port, CI => 
                           SUMB_24_1_port, CO => CARRYB_25_0_port, S => 
                           PRODUCT(25));
   S2_25_1 : FA_X1 port map( A => ab_25_1_port, B => CARRYB_24_1_port, CI => 
                           SUMB_24_2_port, CO => CARRYB_25_1_port, S => 
                           SUMB_25_1_port);
   S2_25_2 : FA_X1 port map( A => ab_25_2_port, B => CARRYB_24_2_port, CI => 
                           SUMB_24_3_port, CO => CARRYB_25_2_port, S => 
                           SUMB_25_2_port);
   S2_25_3 : FA_X1 port map( A => ab_25_3_port, B => CARRYB_24_3_port, CI => 
                           SUMB_24_4_port, CO => CARRYB_25_3_port, S => 
                           SUMB_25_3_port);
   S2_25_4 : FA_X1 port map( A => ab_25_4_port, B => CARRYB_24_4_port, CI => 
                           SUMB_24_5_port, CO => CARRYB_25_4_port, S => 
                           SUMB_25_4_port);
   S2_25_5 : FA_X1 port map( A => ab_25_5_port, B => CARRYB_24_5_port, CI => 
                           SUMB_24_6_port, CO => CARRYB_25_5_port, S => 
                           SUMB_25_5_port);
   S2_25_6 : FA_X1 port map( A => ab_25_6_port, B => CARRYB_24_6_port, CI => 
                           SUMB_24_7_port, CO => n_1039, S => SUMB_25_6_port);
   S1_24_0 : FA_X1 port map( A => ab_24_0_port, B => CARRYB_23_0_port, CI => 
                           SUMB_23_1_port, CO => CARRYB_24_0_port, S => 
                           PRODUCT(24));
   S2_24_1 : FA_X1 port map( A => ab_24_1_port, B => CARRYB_23_1_port, CI => 
                           SUMB_23_2_port, CO => CARRYB_24_1_port, S => 
                           SUMB_24_1_port);
   S2_24_2 : FA_X1 port map( A => ab_24_2_port, B => CARRYB_23_2_port, CI => 
                           SUMB_23_3_port, CO => CARRYB_24_2_port, S => 
                           SUMB_24_2_port);
   S2_24_3 : FA_X1 port map( A => ab_24_3_port, B => CARRYB_23_3_port, CI => 
                           SUMB_23_4_port, CO => CARRYB_24_3_port, S => 
                           SUMB_24_3_port);
   S2_24_4 : FA_X1 port map( A => ab_24_4_port, B => CARRYB_23_4_port, CI => 
                           SUMB_23_5_port, CO => CARRYB_24_4_port, S => 
                           SUMB_24_4_port);
   S2_24_5 : FA_X1 port map( A => ab_24_5_port, B => CARRYB_23_5_port, CI => 
                           SUMB_23_6_port, CO => CARRYB_24_5_port, S => 
                           SUMB_24_5_port);
   S2_24_6 : FA_X1 port map( A => ab_24_6_port, B => CARRYB_23_6_port, CI => 
                           SUMB_23_7_port, CO => CARRYB_24_6_port, S => 
                           SUMB_24_6_port);
   S2_24_7 : FA_X1 port map( A => ab_24_7_port, B => CARRYB_23_7_port, CI => 
                           SUMB_23_8_port, CO => n_1040, S => SUMB_24_7_port);
   S1_23_0 : FA_X1 port map( A => ab_23_0_port, B => CARRYB_22_0_port, CI => 
                           SUMB_22_1_port, CO => CARRYB_23_0_port, S => 
                           PRODUCT(23));
   S2_23_1 : FA_X1 port map( A => ab_23_1_port, B => CARRYB_22_1_port, CI => 
                           SUMB_22_2_port, CO => CARRYB_23_1_port, S => 
                           SUMB_23_1_port);
   S2_23_2 : FA_X1 port map( A => ab_23_2_port, B => CARRYB_22_2_port, CI => 
                           SUMB_22_3_port, CO => CARRYB_23_2_port, S => 
                           SUMB_23_2_port);
   S2_23_3 : FA_X1 port map( A => ab_23_3_port, B => CARRYB_22_3_port, CI => 
                           SUMB_22_4_port, CO => CARRYB_23_3_port, S => 
                           SUMB_23_3_port);
   S2_23_4 : FA_X1 port map( A => ab_23_4_port, B => CARRYB_22_4_port, CI => 
                           SUMB_22_5_port, CO => CARRYB_23_4_port, S => 
                           SUMB_23_4_port);
   S2_23_5 : FA_X1 port map( A => ab_23_5_port, B => CARRYB_22_5_port, CI => 
                           SUMB_22_6_port, CO => CARRYB_23_5_port, S => 
                           SUMB_23_5_port);
   S2_23_6 : FA_X1 port map( A => ab_23_6_port, B => CARRYB_22_6_port, CI => 
                           SUMB_22_7_port, CO => CARRYB_23_6_port, S => 
                           SUMB_23_6_port);
   S2_23_7 : FA_X1 port map( A => ab_23_7_port, B => CARRYB_22_7_port, CI => 
                           SUMB_22_8_port, CO => CARRYB_23_7_port, S => 
                           SUMB_23_7_port);
   S2_23_8 : FA_X1 port map( A => ab_23_8_port, B => CARRYB_22_8_port, CI => 
                           SUMB_22_9_port, CO => n_1041, S => SUMB_23_8_port);
   S1_22_0 : FA_X1 port map( A => ab_22_0_port, B => CARRYB_21_0_port, CI => 
                           SUMB_21_1_port, CO => CARRYB_22_0_port, S => 
                           PRODUCT(22));
   S2_22_1 : FA_X1 port map( A => ab_22_1_port, B => CARRYB_21_1_port, CI => 
                           SUMB_21_2_port, CO => CARRYB_22_1_port, S => 
                           SUMB_22_1_port);
   S2_22_2 : FA_X1 port map( A => ab_22_2_port, B => CARRYB_21_2_port, CI => 
                           SUMB_21_3_port, CO => CARRYB_22_2_port, S => 
                           SUMB_22_2_port);
   S2_22_3 : FA_X1 port map( A => ab_22_3_port, B => CARRYB_21_3_port, CI => 
                           SUMB_21_4_port, CO => CARRYB_22_3_port, S => 
                           SUMB_22_3_port);
   S2_22_4 : FA_X1 port map( A => ab_22_4_port, B => CARRYB_21_4_port, CI => 
                           SUMB_21_5_port, CO => CARRYB_22_4_port, S => 
                           SUMB_22_4_port);
   S2_22_5 : FA_X1 port map( A => ab_22_5_port, B => CARRYB_21_5_port, CI => 
                           SUMB_21_6_port, CO => CARRYB_22_5_port, S => 
                           SUMB_22_5_port);
   S2_22_6 : FA_X1 port map( A => ab_22_6_port, B => CARRYB_21_6_port, CI => 
                           SUMB_21_7_port, CO => CARRYB_22_6_port, S => 
                           SUMB_22_6_port);
   S2_22_7 : FA_X1 port map( A => ab_22_7_port, B => CARRYB_21_7_port, CI => 
                           SUMB_21_8_port, CO => CARRYB_22_7_port, S => 
                           SUMB_22_7_port);
   S2_22_8 : FA_X1 port map( A => ab_22_8_port, B => CARRYB_21_8_port, CI => 
                           SUMB_21_9_port, CO => CARRYB_22_8_port, S => 
                           SUMB_22_8_port);
   S2_22_9 : FA_X1 port map( A => ab_22_9_port, B => CARRYB_21_9_port, CI => 
                           SUMB_21_10_port, CO => n_1042, S => SUMB_22_9_port);
   S1_21_0 : FA_X1 port map( A => ab_21_0_port, B => CARRYB_20_0_port, CI => 
                           SUMB_20_1_port, CO => CARRYB_21_0_port, S => 
                           PRODUCT(21));
   S2_21_1 : FA_X1 port map( A => ab_21_1_port, B => CARRYB_20_1_port, CI => 
                           SUMB_20_2_port, CO => CARRYB_21_1_port, S => 
                           SUMB_21_1_port);
   S2_21_2 : FA_X1 port map( A => ab_21_2_port, B => CARRYB_20_2_port, CI => 
                           SUMB_20_3_port, CO => CARRYB_21_2_port, S => 
                           SUMB_21_2_port);
   S2_21_3 : FA_X1 port map( A => ab_21_3_port, B => CARRYB_20_3_port, CI => 
                           SUMB_20_4_port, CO => CARRYB_21_3_port, S => 
                           SUMB_21_3_port);
   S2_21_4 : FA_X1 port map( A => ab_21_4_port, B => CARRYB_20_4_port, CI => 
                           SUMB_20_5_port, CO => CARRYB_21_4_port, S => 
                           SUMB_21_4_port);
   S2_21_5 : FA_X1 port map( A => ab_21_5_port, B => CARRYB_20_5_port, CI => 
                           SUMB_20_6_port, CO => CARRYB_21_5_port, S => 
                           SUMB_21_5_port);
   S2_21_6 : FA_X1 port map( A => ab_21_6_port, B => CARRYB_20_6_port, CI => 
                           SUMB_20_7_port, CO => CARRYB_21_6_port, S => 
                           SUMB_21_6_port);
   S2_21_7 : FA_X1 port map( A => ab_21_7_port, B => CARRYB_20_7_port, CI => 
                           SUMB_20_8_port, CO => CARRYB_21_7_port, S => 
                           SUMB_21_7_port);
   S2_21_8 : FA_X1 port map( A => ab_21_8_port, B => CARRYB_20_8_port, CI => 
                           SUMB_20_9_port, CO => CARRYB_21_8_port, S => 
                           SUMB_21_8_port);
   S2_21_9 : FA_X1 port map( A => ab_21_9_port, B => CARRYB_20_9_port, CI => 
                           SUMB_20_10_port, CO => CARRYB_21_9_port, S => 
                           SUMB_21_9_port);
   S2_21_10 : FA_X1 port map( A => ab_21_10_port, B => CARRYB_20_10_port, CI =>
                           SUMB_20_11_port, CO => n_1043, S => SUMB_21_10_port)
                           ;
   S1_20_0 : FA_X1 port map( A => ab_20_0_port, B => CARRYB_19_0_port, CI => 
                           SUMB_19_1_port, CO => CARRYB_20_0_port, S => 
                           PRODUCT(20));
   S2_20_1 : FA_X1 port map( A => ab_20_1_port, B => CARRYB_19_1_port, CI => 
                           SUMB_19_2_port, CO => CARRYB_20_1_port, S => 
                           SUMB_20_1_port);
   S2_20_2 : FA_X1 port map( A => ab_20_2_port, B => CARRYB_19_2_port, CI => 
                           SUMB_19_3_port, CO => CARRYB_20_2_port, S => 
                           SUMB_20_2_port);
   S2_20_3 : FA_X1 port map( A => ab_20_3_port, B => CARRYB_19_3_port, CI => 
                           SUMB_19_4_port, CO => CARRYB_20_3_port, S => 
                           SUMB_20_3_port);
   S2_20_4 : FA_X1 port map( A => ab_20_4_port, B => CARRYB_19_4_port, CI => 
                           SUMB_19_5_port, CO => CARRYB_20_4_port, S => 
                           SUMB_20_4_port);
   S2_20_5 : FA_X1 port map( A => ab_20_5_port, B => CARRYB_19_5_port, CI => 
                           SUMB_19_6_port, CO => CARRYB_20_5_port, S => 
                           SUMB_20_5_port);
   S2_20_6 : FA_X1 port map( A => ab_20_6_port, B => CARRYB_19_6_port, CI => 
                           SUMB_19_7_port, CO => CARRYB_20_6_port, S => 
                           SUMB_20_6_port);
   S2_20_7 : FA_X1 port map( A => ab_20_7_port, B => CARRYB_19_7_port, CI => 
                           SUMB_19_8_port, CO => CARRYB_20_7_port, S => 
                           SUMB_20_7_port);
   S2_20_8 : FA_X1 port map( A => ab_20_8_port, B => CARRYB_19_8_port, CI => 
                           SUMB_19_9_port, CO => CARRYB_20_8_port, S => 
                           SUMB_20_8_port);
   S2_20_9 : FA_X1 port map( A => ab_20_9_port, B => CARRYB_19_9_port, CI => 
                           SUMB_19_10_port, CO => CARRYB_20_9_port, S => 
                           SUMB_20_9_port);
   S2_20_10 : FA_X1 port map( A => ab_20_10_port, B => CARRYB_19_10_port, CI =>
                           SUMB_19_11_port, CO => CARRYB_20_10_port, S => 
                           SUMB_20_10_port);
   S2_20_11 : FA_X1 port map( A => ab_20_11_port, B => CARRYB_19_11_port, CI =>
                           SUMB_19_12_port, CO => n_1044, S => SUMB_20_11_port)
                           ;
   S1_19_0 : FA_X1 port map( A => ab_19_0_port, B => CARRYB_18_0_port, CI => 
                           SUMB_18_1_port, CO => CARRYB_19_0_port, S => 
                           PRODUCT(19));
   S2_19_1 : FA_X1 port map( A => ab_19_1_port, B => CARRYB_18_1_port, CI => 
                           SUMB_18_2_port, CO => CARRYB_19_1_port, S => 
                           SUMB_19_1_port);
   S2_19_2 : FA_X1 port map( A => ab_19_2_port, B => CARRYB_18_2_port, CI => 
                           SUMB_18_3_port, CO => CARRYB_19_2_port, S => 
                           SUMB_19_2_port);
   S2_19_3 : FA_X1 port map( A => ab_19_3_port, B => CARRYB_18_3_port, CI => 
                           SUMB_18_4_port, CO => CARRYB_19_3_port, S => 
                           SUMB_19_3_port);
   S2_19_4 : FA_X1 port map( A => ab_19_4_port, B => CARRYB_18_4_port, CI => 
                           SUMB_18_5_port, CO => CARRYB_19_4_port, S => 
                           SUMB_19_4_port);
   S2_19_5 : FA_X1 port map( A => ab_19_5_port, B => CARRYB_18_5_port, CI => 
                           SUMB_18_6_port, CO => CARRYB_19_5_port, S => 
                           SUMB_19_5_port);
   S2_19_6 : FA_X1 port map( A => ab_19_6_port, B => CARRYB_18_6_port, CI => 
                           SUMB_18_7_port, CO => CARRYB_19_6_port, S => 
                           SUMB_19_6_port);
   S2_19_7 : FA_X1 port map( A => ab_19_7_port, B => CARRYB_18_7_port, CI => 
                           SUMB_18_8_port, CO => CARRYB_19_7_port, S => 
                           SUMB_19_7_port);
   S2_19_8 : FA_X1 port map( A => ab_19_8_port, B => CARRYB_18_8_port, CI => 
                           SUMB_18_9_port, CO => CARRYB_19_8_port, S => 
                           SUMB_19_8_port);
   S2_19_9 : FA_X1 port map( A => ab_19_9_port, B => CARRYB_18_9_port, CI => 
                           SUMB_18_10_port, CO => CARRYB_19_9_port, S => 
                           SUMB_19_9_port);
   S2_19_10 : FA_X1 port map( A => ab_19_10_port, B => CARRYB_18_10_port, CI =>
                           SUMB_18_11_port, CO => CARRYB_19_10_port, S => 
                           SUMB_19_10_port);
   S2_19_11 : FA_X1 port map( A => ab_19_11_port, B => CARRYB_18_11_port, CI =>
                           SUMB_18_12_port, CO => CARRYB_19_11_port, S => 
                           SUMB_19_11_port);
   S2_19_12 : FA_X1 port map( A => ab_19_12_port, B => CARRYB_18_12_port, CI =>
                           SUMB_18_13_port, CO => n_1045, S => SUMB_19_12_port)
                           ;
   S1_18_0 : FA_X1 port map( A => ab_18_0_port, B => CARRYB_17_0_port, CI => 
                           SUMB_17_1_port, CO => CARRYB_18_0_port, S => 
                           PRODUCT(18));
   S2_18_1 : FA_X1 port map( A => ab_18_1_port, B => CARRYB_17_1_port, CI => 
                           SUMB_17_2_port, CO => CARRYB_18_1_port, S => 
                           SUMB_18_1_port);
   S2_18_2 : FA_X1 port map( A => ab_18_2_port, B => CARRYB_17_2_port, CI => 
                           SUMB_17_3_port, CO => CARRYB_18_2_port, S => 
                           SUMB_18_2_port);
   S2_18_3 : FA_X1 port map( A => ab_18_3_port, B => CARRYB_17_3_port, CI => 
                           SUMB_17_4_port, CO => CARRYB_18_3_port, S => 
                           SUMB_18_3_port);
   S2_18_4 : FA_X1 port map( A => ab_18_4_port, B => CARRYB_17_4_port, CI => 
                           SUMB_17_5_port, CO => CARRYB_18_4_port, S => 
                           SUMB_18_4_port);
   S2_18_5 : FA_X1 port map( A => ab_18_5_port, B => CARRYB_17_5_port, CI => 
                           SUMB_17_6_port, CO => CARRYB_18_5_port, S => 
                           SUMB_18_5_port);
   S2_18_6 : FA_X1 port map( A => ab_18_6_port, B => CARRYB_17_6_port, CI => 
                           SUMB_17_7_port, CO => CARRYB_18_6_port, S => 
                           SUMB_18_6_port);
   S2_18_7 : FA_X1 port map( A => ab_18_7_port, B => CARRYB_17_7_port, CI => 
                           SUMB_17_8_port, CO => CARRYB_18_7_port, S => 
                           SUMB_18_7_port);
   S2_18_8 : FA_X1 port map( A => ab_18_8_port, B => CARRYB_17_8_port, CI => 
                           SUMB_17_9_port, CO => CARRYB_18_8_port, S => 
                           SUMB_18_8_port);
   S2_18_9 : FA_X1 port map( A => ab_18_9_port, B => CARRYB_17_9_port, CI => 
                           SUMB_17_10_port, CO => CARRYB_18_9_port, S => 
                           SUMB_18_9_port);
   S2_18_10 : FA_X1 port map( A => ab_18_10_port, B => CARRYB_17_10_port, CI =>
                           SUMB_17_11_port, CO => CARRYB_18_10_port, S => 
                           SUMB_18_10_port);
   S2_18_11 : FA_X1 port map( A => ab_18_11_port, B => CARRYB_17_11_port, CI =>
                           SUMB_17_12_port, CO => CARRYB_18_11_port, S => 
                           SUMB_18_11_port);
   S2_18_12 : FA_X1 port map( A => ab_18_12_port, B => CARRYB_17_12_port, CI =>
                           SUMB_17_13_port, CO => CARRYB_18_12_port, S => 
                           SUMB_18_12_port);
   S2_18_13 : FA_X1 port map( A => ab_18_13_port, B => CARRYB_17_13_port, CI =>
                           SUMB_17_14_port, CO => n_1046, S => SUMB_18_13_port)
                           ;
   S1_17_0 : FA_X1 port map( A => ab_17_0_port, B => CARRYB_16_0_port, CI => 
                           SUMB_16_1_port, CO => CARRYB_17_0_port, S => 
                           PRODUCT(17));
   S2_17_1 : FA_X1 port map( A => ab_17_1_port, B => CARRYB_16_1_port, CI => 
                           SUMB_16_2_port, CO => CARRYB_17_1_port, S => 
                           SUMB_17_1_port);
   S2_17_2 : FA_X1 port map( A => ab_17_2_port, B => CARRYB_16_2_port, CI => 
                           SUMB_16_3_port, CO => CARRYB_17_2_port, S => 
                           SUMB_17_2_port);
   S2_17_3 : FA_X1 port map( A => ab_17_3_port, B => CARRYB_16_3_port, CI => 
                           SUMB_16_4_port, CO => CARRYB_17_3_port, S => 
                           SUMB_17_3_port);
   S2_17_4 : FA_X1 port map( A => ab_17_4_port, B => CARRYB_16_4_port, CI => 
                           SUMB_16_5_port, CO => CARRYB_17_4_port, S => 
                           SUMB_17_4_port);
   S2_17_5 : FA_X1 port map( A => ab_17_5_port, B => CARRYB_16_5_port, CI => 
                           SUMB_16_6_port, CO => CARRYB_17_5_port, S => 
                           SUMB_17_5_port);
   S2_17_6 : FA_X1 port map( A => ab_17_6_port, B => CARRYB_16_6_port, CI => 
                           SUMB_16_7_port, CO => CARRYB_17_6_port, S => 
                           SUMB_17_6_port);
   S2_17_7 : FA_X1 port map( A => ab_17_7_port, B => CARRYB_16_7_port, CI => 
                           SUMB_16_8_port, CO => CARRYB_17_7_port, S => 
                           SUMB_17_7_port);
   S2_17_8 : FA_X1 port map( A => ab_17_8_port, B => CARRYB_16_8_port, CI => 
                           SUMB_16_9_port, CO => CARRYB_17_8_port, S => 
                           SUMB_17_8_port);
   S2_17_9 : FA_X1 port map( A => ab_17_9_port, B => CARRYB_16_9_port, CI => 
                           SUMB_16_10_port, CO => CARRYB_17_9_port, S => 
                           SUMB_17_9_port);
   S2_17_10 : FA_X1 port map( A => ab_17_10_port, B => CARRYB_16_10_port, CI =>
                           SUMB_16_11_port, CO => CARRYB_17_10_port, S => 
                           SUMB_17_10_port);
   S2_17_11 : FA_X1 port map( A => ab_17_11_port, B => CARRYB_16_11_port, CI =>
                           SUMB_16_12_port, CO => CARRYB_17_11_port, S => 
                           SUMB_17_11_port);
   S2_17_12 : FA_X1 port map( A => ab_17_12_port, B => CARRYB_16_12_port, CI =>
                           SUMB_16_13_port, CO => CARRYB_17_12_port, S => 
                           SUMB_17_12_port);
   S2_17_13 : FA_X1 port map( A => ab_17_13_port, B => CARRYB_16_13_port, CI =>
                           SUMB_16_14_port, CO => CARRYB_17_13_port, S => 
                           SUMB_17_13_port);
   S2_17_14 : FA_X1 port map( A => ab_17_14_port, B => CARRYB_16_14_port, CI =>
                           SUMB_16_15_port, CO => n_1047, S => SUMB_17_14_port)
                           ;
   S1_16_0 : FA_X1 port map( A => ab_16_0_port, B => CARRYB_15_0_port, CI => 
                           SUMB_15_1_port, CO => CARRYB_16_0_port, S => 
                           PRODUCT(16));
   S2_16_1 : FA_X1 port map( A => ab_16_1_port, B => CARRYB_15_1_port, CI => 
                           SUMB_15_2_port, CO => CARRYB_16_1_port, S => 
                           SUMB_16_1_port);
   S2_16_2 : FA_X1 port map( A => ab_16_2_port, B => CARRYB_15_2_port, CI => 
                           SUMB_15_3_port, CO => CARRYB_16_2_port, S => 
                           SUMB_16_2_port);
   S2_16_3 : FA_X1 port map( A => ab_16_3_port, B => CARRYB_15_3_port, CI => 
                           SUMB_15_4_port, CO => CARRYB_16_3_port, S => 
                           SUMB_16_3_port);
   S2_16_4 : FA_X1 port map( A => ab_16_4_port, B => CARRYB_15_4_port, CI => 
                           SUMB_15_5_port, CO => CARRYB_16_4_port, S => 
                           SUMB_16_4_port);
   S2_16_5 : FA_X1 port map( A => ab_16_5_port, B => CARRYB_15_5_port, CI => 
                           SUMB_15_6_port, CO => CARRYB_16_5_port, S => 
                           SUMB_16_5_port);
   S2_16_6 : FA_X1 port map( A => ab_16_6_port, B => CARRYB_15_6_port, CI => 
                           SUMB_15_7_port, CO => CARRYB_16_6_port, S => 
                           SUMB_16_6_port);
   S2_16_7 : FA_X1 port map( A => ab_16_7_port, B => CARRYB_15_7_port, CI => 
                           SUMB_15_8_port, CO => CARRYB_16_7_port, S => 
                           SUMB_16_7_port);
   S2_16_8 : FA_X1 port map( A => ab_16_8_port, B => CARRYB_15_8_port, CI => 
                           SUMB_15_9_port, CO => CARRYB_16_8_port, S => 
                           SUMB_16_8_port);
   S2_16_9 : FA_X1 port map( A => ab_16_9_port, B => CARRYB_15_9_port, CI => 
                           SUMB_15_10_port, CO => CARRYB_16_9_port, S => 
                           SUMB_16_9_port);
   S2_16_10 : FA_X1 port map( A => ab_16_10_port, B => CARRYB_15_10_port, CI =>
                           SUMB_15_11_port, CO => CARRYB_16_10_port, S => 
                           SUMB_16_10_port);
   S2_16_11 : FA_X1 port map( A => ab_16_11_port, B => CARRYB_15_11_port, CI =>
                           SUMB_15_12_port, CO => CARRYB_16_11_port, S => 
                           SUMB_16_11_port);
   S2_16_12 : FA_X1 port map( A => ab_16_12_port, B => CARRYB_15_12_port, CI =>
                           SUMB_15_13_port, CO => CARRYB_16_12_port, S => 
                           SUMB_16_12_port);
   S2_16_13 : FA_X1 port map( A => ab_16_13_port, B => CARRYB_15_13_port, CI =>
                           SUMB_15_14_port, CO => CARRYB_16_13_port, S => 
                           SUMB_16_13_port);
   S2_16_14 : FA_X1 port map( A => ab_16_14_port, B => CARRYB_15_14_port, CI =>
                           SUMB_15_15_port, CO => CARRYB_16_14_port, S => 
                           SUMB_16_14_port);
   S2_16_15 : FA_X1 port map( A => ab_16_15_port, B => CARRYB_15_15_port, CI =>
                           SUMB_15_16_port, CO => n_1048, S => SUMB_16_15_port)
                           ;
   S1_15_0 : FA_X1 port map( A => ab_15_0_port, B => CARRYB_14_0_port, CI => 
                           SUMB_14_1_port, CO => CARRYB_15_0_port, S => 
                           PRODUCT(15));
   S2_15_1 : FA_X1 port map( A => ab_15_1_port, B => CARRYB_14_1_port, CI => 
                           SUMB_14_2_port, CO => CARRYB_15_1_port, S => 
                           SUMB_15_1_port);
   S2_15_2 : FA_X1 port map( A => ab_15_2_port, B => CARRYB_14_2_port, CI => 
                           SUMB_14_3_port, CO => CARRYB_15_2_port, S => 
                           SUMB_15_2_port);
   S2_15_3 : FA_X1 port map( A => ab_15_3_port, B => CARRYB_14_3_port, CI => 
                           SUMB_14_4_port, CO => CARRYB_15_3_port, S => 
                           SUMB_15_3_port);
   S2_15_4 : FA_X1 port map( A => ab_15_4_port, B => CARRYB_14_4_port, CI => 
                           SUMB_14_5_port, CO => CARRYB_15_4_port, S => 
                           SUMB_15_4_port);
   S2_15_5 : FA_X1 port map( A => ab_15_5_port, B => CARRYB_14_5_port, CI => 
                           SUMB_14_6_port, CO => CARRYB_15_5_port, S => 
                           SUMB_15_5_port);
   S2_15_6 : FA_X1 port map( A => ab_15_6_port, B => CARRYB_14_6_port, CI => 
                           SUMB_14_7_port, CO => CARRYB_15_6_port, S => 
                           SUMB_15_6_port);
   S2_15_7 : FA_X1 port map( A => ab_15_7_port, B => CARRYB_14_7_port, CI => 
                           SUMB_14_8_port, CO => CARRYB_15_7_port, S => 
                           SUMB_15_7_port);
   S2_15_8 : FA_X1 port map( A => ab_15_8_port, B => CARRYB_14_8_port, CI => 
                           SUMB_14_9_port, CO => CARRYB_15_8_port, S => 
                           SUMB_15_8_port);
   S2_15_9 : FA_X1 port map( A => ab_15_9_port, B => CARRYB_14_9_port, CI => 
                           SUMB_14_10_port, CO => CARRYB_15_9_port, S => 
                           SUMB_15_9_port);
   S2_15_10 : FA_X1 port map( A => ab_15_10_port, B => CARRYB_14_10_port, CI =>
                           SUMB_14_11_port, CO => CARRYB_15_10_port, S => 
                           SUMB_15_10_port);
   S2_15_11 : FA_X1 port map( A => ab_15_11_port, B => CARRYB_14_11_port, CI =>
                           SUMB_14_12_port, CO => CARRYB_15_11_port, S => 
                           SUMB_15_11_port);
   S2_15_12 : FA_X1 port map( A => ab_15_12_port, B => CARRYB_14_12_port, CI =>
                           SUMB_14_13_port, CO => CARRYB_15_12_port, S => 
                           SUMB_15_12_port);
   S2_15_13 : FA_X1 port map( A => ab_15_13_port, B => CARRYB_14_13_port, CI =>
                           SUMB_14_14_port, CO => CARRYB_15_13_port, S => 
                           SUMB_15_13_port);
   S2_15_14 : FA_X1 port map( A => ab_15_14_port, B => CARRYB_14_14_port, CI =>
                           SUMB_14_15_port, CO => CARRYB_15_14_port, S => 
                           SUMB_15_14_port);
   S2_15_15 : FA_X1 port map( A => ab_15_15_port, B => CARRYB_14_15_port, CI =>
                           SUMB_14_16_port, CO => CARRYB_15_15_port, S => 
                           SUMB_15_15_port);
   S2_15_16 : FA_X1 port map( A => ab_15_16_port, B => CARRYB_14_16_port, CI =>
                           SUMB_14_17_port, CO => n_1049, S => SUMB_15_16_port)
                           ;
   S1_14_0 : FA_X1 port map( A => ab_14_0_port, B => CARRYB_13_0_port, CI => 
                           SUMB_13_1_port, CO => CARRYB_14_0_port, S => 
                           PRODUCT(14));
   S2_14_1 : FA_X1 port map( A => ab_14_1_port, B => CARRYB_13_1_port, CI => 
                           SUMB_13_2_port, CO => CARRYB_14_1_port, S => 
                           SUMB_14_1_port);
   S2_14_2 : FA_X1 port map( A => ab_14_2_port, B => CARRYB_13_2_port, CI => 
                           SUMB_13_3_port, CO => CARRYB_14_2_port, S => 
                           SUMB_14_2_port);
   S2_14_3 : FA_X1 port map( A => ab_14_3_port, B => CARRYB_13_3_port, CI => 
                           SUMB_13_4_port, CO => CARRYB_14_3_port, S => 
                           SUMB_14_3_port);
   S2_14_4 : FA_X1 port map( A => ab_14_4_port, B => CARRYB_13_4_port, CI => 
                           SUMB_13_5_port, CO => CARRYB_14_4_port, S => 
                           SUMB_14_4_port);
   S2_14_5 : FA_X1 port map( A => ab_14_5_port, B => CARRYB_13_5_port, CI => 
                           SUMB_13_6_port, CO => CARRYB_14_5_port, S => 
                           SUMB_14_5_port);
   S2_14_6 : FA_X1 port map( A => ab_14_6_port, B => CARRYB_13_6_port, CI => 
                           SUMB_13_7_port, CO => CARRYB_14_6_port, S => 
                           SUMB_14_6_port);
   S2_14_7 : FA_X1 port map( A => ab_14_7_port, B => CARRYB_13_7_port, CI => 
                           SUMB_13_8_port, CO => CARRYB_14_7_port, S => 
                           SUMB_14_7_port);
   S2_14_8 : FA_X1 port map( A => ab_14_8_port, B => CARRYB_13_8_port, CI => 
                           SUMB_13_9_port, CO => CARRYB_14_8_port, S => 
                           SUMB_14_8_port);
   S2_14_9 : FA_X1 port map( A => ab_14_9_port, B => CARRYB_13_9_port, CI => 
                           SUMB_13_10_port, CO => CARRYB_14_9_port, S => 
                           SUMB_14_9_port);
   S2_14_10 : FA_X1 port map( A => ab_14_10_port, B => CARRYB_13_10_port, CI =>
                           SUMB_13_11_port, CO => CARRYB_14_10_port, S => 
                           SUMB_14_10_port);
   S2_14_11 : FA_X1 port map( A => ab_14_11_port, B => CARRYB_13_11_port, CI =>
                           SUMB_13_12_port, CO => CARRYB_14_11_port, S => 
                           SUMB_14_11_port);
   S2_14_12 : FA_X1 port map( A => ab_14_12_port, B => CARRYB_13_12_port, CI =>
                           SUMB_13_13_port, CO => CARRYB_14_12_port, S => 
                           SUMB_14_12_port);
   S2_14_13 : FA_X1 port map( A => ab_14_13_port, B => CARRYB_13_13_port, CI =>
                           SUMB_13_14_port, CO => CARRYB_14_13_port, S => 
                           SUMB_14_13_port);
   S2_14_14 : FA_X1 port map( A => ab_14_14_port, B => CARRYB_13_14_port, CI =>
                           SUMB_13_15_port, CO => CARRYB_14_14_port, S => 
                           SUMB_14_14_port);
   S2_14_15 : FA_X1 port map( A => ab_14_15_port, B => CARRYB_13_15_port, CI =>
                           SUMB_13_16_port, CO => CARRYB_14_15_port, S => 
                           SUMB_14_15_port);
   S2_14_16 : FA_X1 port map( A => ab_14_16_port, B => CARRYB_13_16_port, CI =>
                           SUMB_13_17_port, CO => CARRYB_14_16_port, S => 
                           SUMB_14_16_port);
   S2_14_17 : FA_X1 port map( A => ab_14_17_port, B => CARRYB_13_17_port, CI =>
                           SUMB_13_18_port, CO => n_1050, S => SUMB_14_17_port)
                           ;
   S1_13_0 : FA_X1 port map( A => ab_13_0_port, B => CARRYB_12_0_port, CI => 
                           SUMB_12_1_port, CO => CARRYB_13_0_port, S => 
                           PRODUCT(13));
   S2_13_1 : FA_X1 port map( A => ab_13_1_port, B => CARRYB_12_1_port, CI => 
                           SUMB_12_2_port, CO => CARRYB_13_1_port, S => 
                           SUMB_13_1_port);
   S2_13_2 : FA_X1 port map( A => ab_13_2_port, B => CARRYB_12_2_port, CI => 
                           SUMB_12_3_port, CO => CARRYB_13_2_port, S => 
                           SUMB_13_2_port);
   S2_13_3 : FA_X1 port map( A => ab_13_3_port, B => CARRYB_12_3_port, CI => 
                           SUMB_12_4_port, CO => CARRYB_13_3_port, S => 
                           SUMB_13_3_port);
   S2_13_4 : FA_X1 port map( A => ab_13_4_port, B => CARRYB_12_4_port, CI => 
                           SUMB_12_5_port, CO => CARRYB_13_4_port, S => 
                           SUMB_13_4_port);
   S2_13_5 : FA_X1 port map( A => ab_13_5_port, B => CARRYB_12_5_port, CI => 
                           SUMB_12_6_port, CO => CARRYB_13_5_port, S => 
                           SUMB_13_5_port);
   S2_13_6 : FA_X1 port map( A => ab_13_6_port, B => CARRYB_12_6_port, CI => 
                           SUMB_12_7_port, CO => CARRYB_13_6_port, S => 
                           SUMB_13_6_port);
   S2_13_7 : FA_X1 port map( A => ab_13_7_port, B => CARRYB_12_7_port, CI => 
                           SUMB_12_8_port, CO => CARRYB_13_7_port, S => 
                           SUMB_13_7_port);
   S2_13_8 : FA_X1 port map( A => ab_13_8_port, B => CARRYB_12_8_port, CI => 
                           SUMB_12_9_port, CO => CARRYB_13_8_port, S => 
                           SUMB_13_8_port);
   S2_13_9 : FA_X1 port map( A => ab_13_9_port, B => CARRYB_12_9_port, CI => 
                           SUMB_12_10_port, CO => CARRYB_13_9_port, S => 
                           SUMB_13_9_port);
   S2_13_10 : FA_X1 port map( A => ab_13_10_port, B => CARRYB_12_10_port, CI =>
                           SUMB_12_11_port, CO => CARRYB_13_10_port, S => 
                           SUMB_13_10_port);
   S2_13_11 : FA_X1 port map( A => ab_13_11_port, B => CARRYB_12_11_port, CI =>
                           SUMB_12_12_port, CO => CARRYB_13_11_port, S => 
                           SUMB_13_11_port);
   S2_13_12 : FA_X1 port map( A => ab_13_12_port, B => CARRYB_12_12_port, CI =>
                           SUMB_12_13_port, CO => CARRYB_13_12_port, S => 
                           SUMB_13_12_port);
   S2_13_13 : FA_X1 port map( A => ab_13_13_port, B => CARRYB_12_13_port, CI =>
                           SUMB_12_14_port, CO => CARRYB_13_13_port, S => 
                           SUMB_13_13_port);
   S2_13_14 : FA_X1 port map( A => ab_13_14_port, B => CARRYB_12_14_port, CI =>
                           SUMB_12_15_port, CO => CARRYB_13_14_port, S => 
                           SUMB_13_14_port);
   S2_13_15 : FA_X1 port map( A => ab_13_15_port, B => CARRYB_12_15_port, CI =>
                           SUMB_12_16_port, CO => CARRYB_13_15_port, S => 
                           SUMB_13_15_port);
   S2_13_16 : FA_X1 port map( A => ab_13_16_port, B => CARRYB_12_16_port, CI =>
                           SUMB_12_17_port, CO => CARRYB_13_16_port, S => 
                           SUMB_13_16_port);
   S2_13_17 : FA_X1 port map( A => ab_13_17_port, B => CARRYB_12_17_port, CI =>
                           SUMB_12_18_port, CO => CARRYB_13_17_port, S => 
                           SUMB_13_17_port);
   S2_13_18 : FA_X1 port map( A => ab_13_18_port, B => CARRYB_12_18_port, CI =>
                           SUMB_12_19_port, CO => n_1051, S => SUMB_13_18_port)
                           ;
   S1_12_0 : FA_X1 port map( A => ab_12_0_port, B => CARRYB_11_0_port, CI => 
                           SUMB_11_1_port, CO => CARRYB_12_0_port, S => 
                           PRODUCT(12));
   S2_12_1 : FA_X1 port map( A => ab_12_1_port, B => CARRYB_11_1_port, CI => 
                           SUMB_11_2_port, CO => CARRYB_12_1_port, S => 
                           SUMB_12_1_port);
   S2_12_2 : FA_X1 port map( A => ab_12_2_port, B => CARRYB_11_2_port, CI => 
                           SUMB_11_3_port, CO => CARRYB_12_2_port, S => 
                           SUMB_12_2_port);
   S2_12_3 : FA_X1 port map( A => ab_12_3_port, B => CARRYB_11_3_port, CI => 
                           SUMB_11_4_port, CO => CARRYB_12_3_port, S => 
                           SUMB_12_3_port);
   S2_12_4 : FA_X1 port map( A => ab_12_4_port, B => CARRYB_11_4_port, CI => 
                           SUMB_11_5_port, CO => CARRYB_12_4_port, S => 
                           SUMB_12_4_port);
   S2_12_5 : FA_X1 port map( A => ab_12_5_port, B => CARRYB_11_5_port, CI => 
                           SUMB_11_6_port, CO => CARRYB_12_5_port, S => 
                           SUMB_12_5_port);
   S2_12_6 : FA_X1 port map( A => ab_12_6_port, B => CARRYB_11_6_port, CI => 
                           SUMB_11_7_port, CO => CARRYB_12_6_port, S => 
                           SUMB_12_6_port);
   S2_12_7 : FA_X1 port map( A => ab_12_7_port, B => CARRYB_11_7_port, CI => 
                           SUMB_11_8_port, CO => CARRYB_12_7_port, S => 
                           SUMB_12_7_port);
   S2_12_8 : FA_X1 port map( A => ab_12_8_port, B => CARRYB_11_8_port, CI => 
                           SUMB_11_9_port, CO => CARRYB_12_8_port, S => 
                           SUMB_12_8_port);
   S2_12_9 : FA_X1 port map( A => ab_12_9_port, B => CARRYB_11_9_port, CI => 
                           SUMB_11_10_port, CO => CARRYB_12_9_port, S => 
                           SUMB_12_9_port);
   S2_12_10 : FA_X1 port map( A => ab_12_10_port, B => CARRYB_11_10_port, CI =>
                           SUMB_11_11_port, CO => CARRYB_12_10_port, S => 
                           SUMB_12_10_port);
   S2_12_11 : FA_X1 port map( A => ab_12_11_port, B => CARRYB_11_11_port, CI =>
                           SUMB_11_12_port, CO => CARRYB_12_11_port, S => 
                           SUMB_12_11_port);
   S2_12_12 : FA_X1 port map( A => ab_12_12_port, B => CARRYB_11_12_port, CI =>
                           SUMB_11_13_port, CO => CARRYB_12_12_port, S => 
                           SUMB_12_12_port);
   S2_12_13 : FA_X1 port map( A => ab_12_13_port, B => CARRYB_11_13_port, CI =>
                           SUMB_11_14_port, CO => CARRYB_12_13_port, S => 
                           SUMB_12_13_port);
   S2_12_14 : FA_X1 port map( A => ab_12_14_port, B => CARRYB_11_14_port, CI =>
                           SUMB_11_15_port, CO => CARRYB_12_14_port, S => 
                           SUMB_12_14_port);
   S2_12_15 : FA_X1 port map( A => ab_12_15_port, B => CARRYB_11_15_port, CI =>
                           SUMB_11_16_port, CO => CARRYB_12_15_port, S => 
                           SUMB_12_15_port);
   S2_12_16 : FA_X1 port map( A => ab_12_16_port, B => CARRYB_11_16_port, CI =>
                           SUMB_11_17_port, CO => CARRYB_12_16_port, S => 
                           SUMB_12_16_port);
   S2_12_17 : FA_X1 port map( A => ab_12_17_port, B => CARRYB_11_17_port, CI =>
                           SUMB_11_18_port, CO => CARRYB_12_17_port, S => 
                           SUMB_12_17_port);
   S2_12_18 : FA_X1 port map( A => ab_12_18_port, B => CARRYB_11_18_port, CI =>
                           SUMB_11_19_port, CO => CARRYB_12_18_port, S => 
                           SUMB_12_18_port);
   S2_12_19 : FA_X1 port map( A => ab_12_19_port, B => CARRYB_11_19_port, CI =>
                           SUMB_11_20_port, CO => n_1052, S => SUMB_12_19_port)
                           ;
   S1_11_0 : FA_X1 port map( A => ab_11_0_port, B => CARRYB_10_0_port, CI => 
                           SUMB_10_1_port, CO => CARRYB_11_0_port, S => 
                           PRODUCT(11));
   S2_11_1 : FA_X1 port map( A => ab_11_1_port, B => CARRYB_10_1_port, CI => 
                           SUMB_10_2_port, CO => CARRYB_11_1_port, S => 
                           SUMB_11_1_port);
   S2_11_2 : FA_X1 port map( A => ab_11_2_port, B => CARRYB_10_2_port, CI => 
                           SUMB_10_3_port, CO => CARRYB_11_2_port, S => 
                           SUMB_11_2_port);
   S2_11_3 : FA_X1 port map( A => ab_11_3_port, B => CARRYB_10_3_port, CI => 
                           SUMB_10_4_port, CO => CARRYB_11_3_port, S => 
                           SUMB_11_3_port);
   S2_11_4 : FA_X1 port map( A => ab_11_4_port, B => CARRYB_10_4_port, CI => 
                           SUMB_10_5_port, CO => CARRYB_11_4_port, S => 
                           SUMB_11_4_port);
   S2_11_5 : FA_X1 port map( A => ab_11_5_port, B => CARRYB_10_5_port, CI => 
                           SUMB_10_6_port, CO => CARRYB_11_5_port, S => 
                           SUMB_11_5_port);
   S2_11_6 : FA_X1 port map( A => ab_11_6_port, B => CARRYB_10_6_port, CI => 
                           SUMB_10_7_port, CO => CARRYB_11_6_port, S => 
                           SUMB_11_6_port);
   S2_11_7 : FA_X1 port map( A => ab_11_7_port, B => CARRYB_10_7_port, CI => 
                           SUMB_10_8_port, CO => CARRYB_11_7_port, S => 
                           SUMB_11_7_port);
   S2_11_8 : FA_X1 port map( A => ab_11_8_port, B => CARRYB_10_8_port, CI => 
                           SUMB_10_9_port, CO => CARRYB_11_8_port, S => 
                           SUMB_11_8_port);
   S2_11_9 : FA_X1 port map( A => ab_11_9_port, B => CARRYB_10_9_port, CI => 
                           SUMB_10_10_port, CO => CARRYB_11_9_port, S => 
                           SUMB_11_9_port);
   S2_11_10 : FA_X1 port map( A => ab_11_10_port, B => CARRYB_10_10_port, CI =>
                           SUMB_10_11_port, CO => CARRYB_11_10_port, S => 
                           SUMB_11_10_port);
   S2_11_11 : FA_X1 port map( A => ab_11_11_port, B => CARRYB_10_11_port, CI =>
                           SUMB_10_12_port, CO => CARRYB_11_11_port, S => 
                           SUMB_11_11_port);
   S2_11_12 : FA_X1 port map( A => ab_11_12_port, B => CARRYB_10_12_port, CI =>
                           SUMB_10_13_port, CO => CARRYB_11_12_port, S => 
                           SUMB_11_12_port);
   S2_11_13 : FA_X1 port map( A => ab_11_13_port, B => CARRYB_10_13_port, CI =>
                           SUMB_10_14_port, CO => CARRYB_11_13_port, S => 
                           SUMB_11_13_port);
   S2_11_14 : FA_X1 port map( A => ab_11_14_port, B => CARRYB_10_14_port, CI =>
                           SUMB_10_15_port, CO => CARRYB_11_14_port, S => 
                           SUMB_11_14_port);
   S2_11_15 : FA_X1 port map( A => ab_11_15_port, B => CARRYB_10_15_port, CI =>
                           SUMB_10_16_port, CO => CARRYB_11_15_port, S => 
                           SUMB_11_15_port);
   S2_11_16 : FA_X1 port map( A => ab_11_16_port, B => CARRYB_10_16_port, CI =>
                           SUMB_10_17_port, CO => CARRYB_11_16_port, S => 
                           SUMB_11_16_port);
   S2_11_17 : FA_X1 port map( A => ab_11_17_port, B => CARRYB_10_17_port, CI =>
                           SUMB_10_18_port, CO => CARRYB_11_17_port, S => 
                           SUMB_11_17_port);
   S2_11_18 : FA_X1 port map( A => ab_11_18_port, B => CARRYB_10_18_port, CI =>
                           SUMB_10_19_port, CO => CARRYB_11_18_port, S => 
                           SUMB_11_18_port);
   S2_11_19 : FA_X1 port map( A => ab_11_19_port, B => CARRYB_10_19_port, CI =>
                           SUMB_10_20_port, CO => CARRYB_11_19_port, S => 
                           SUMB_11_19_port);
   S2_11_20 : FA_X1 port map( A => ab_11_20_port, B => CARRYB_10_20_port, CI =>
                           SUMB_10_21_port, CO => n_1053, S => SUMB_11_20_port)
                           ;
   S1_10_0 : FA_X1 port map( A => ab_10_0_port, B => CARRYB_9_0_port, CI => 
                           SUMB_9_1_port, CO => CARRYB_10_0_port, S => 
                           PRODUCT(10));
   S2_10_1 : FA_X1 port map( A => ab_10_1_port, B => CARRYB_9_1_port, CI => 
                           SUMB_9_2_port, CO => CARRYB_10_1_port, S => 
                           SUMB_10_1_port);
   S2_10_2 : FA_X1 port map( A => ab_10_2_port, B => CARRYB_9_2_port, CI => 
                           SUMB_9_3_port, CO => CARRYB_10_2_port, S => 
                           SUMB_10_2_port);
   S2_10_3 : FA_X1 port map( A => ab_10_3_port, B => CARRYB_9_3_port, CI => 
                           SUMB_9_4_port, CO => CARRYB_10_3_port, S => 
                           SUMB_10_3_port);
   S2_10_4 : FA_X1 port map( A => ab_10_4_port, B => CARRYB_9_4_port, CI => 
                           SUMB_9_5_port, CO => CARRYB_10_4_port, S => 
                           SUMB_10_4_port);
   S2_10_5 : FA_X1 port map( A => ab_10_5_port, B => CARRYB_9_5_port, CI => 
                           SUMB_9_6_port, CO => CARRYB_10_5_port, S => 
                           SUMB_10_5_port);
   S2_10_6 : FA_X1 port map( A => ab_10_6_port, B => CARRYB_9_6_port, CI => 
                           SUMB_9_7_port, CO => CARRYB_10_6_port, S => 
                           SUMB_10_6_port);
   S2_10_7 : FA_X1 port map( A => ab_10_7_port, B => CARRYB_9_7_port, CI => 
                           SUMB_9_8_port, CO => CARRYB_10_7_port, S => 
                           SUMB_10_7_port);
   S2_10_8 : FA_X1 port map( A => ab_10_8_port, B => CARRYB_9_8_port, CI => 
                           SUMB_9_9_port, CO => CARRYB_10_8_port, S => 
                           SUMB_10_8_port);
   S2_10_9 : FA_X1 port map( A => ab_10_9_port, B => CARRYB_9_9_port, CI => 
                           SUMB_9_10_port, CO => CARRYB_10_9_port, S => 
                           SUMB_10_9_port);
   S2_10_10 : FA_X1 port map( A => ab_10_10_port, B => CARRYB_9_10_port, CI => 
                           SUMB_9_11_port, CO => CARRYB_10_10_port, S => 
                           SUMB_10_10_port);
   S2_10_11 : FA_X1 port map( A => ab_10_11_port, B => CARRYB_9_11_port, CI => 
                           SUMB_9_12_port, CO => CARRYB_10_11_port, S => 
                           SUMB_10_11_port);
   S2_10_12 : FA_X1 port map( A => ab_10_12_port, B => CARRYB_9_12_port, CI => 
                           SUMB_9_13_port, CO => CARRYB_10_12_port, S => 
                           SUMB_10_12_port);
   S2_10_13 : FA_X1 port map( A => ab_10_13_port, B => CARRYB_9_13_port, CI => 
                           SUMB_9_14_port, CO => CARRYB_10_13_port, S => 
                           SUMB_10_13_port);
   S2_10_14 : FA_X1 port map( A => ab_10_14_port, B => CARRYB_9_14_port, CI => 
                           SUMB_9_15_port, CO => CARRYB_10_14_port, S => 
                           SUMB_10_14_port);
   S2_10_15 : FA_X1 port map( A => ab_10_15_port, B => CARRYB_9_15_port, CI => 
                           SUMB_9_16_port, CO => CARRYB_10_15_port, S => 
                           SUMB_10_15_port);
   S2_10_16 : FA_X1 port map( A => ab_10_16_port, B => CARRYB_9_16_port, CI => 
                           SUMB_9_17_port, CO => CARRYB_10_16_port, S => 
                           SUMB_10_16_port);
   S2_10_17 : FA_X1 port map( A => ab_10_17_port, B => CARRYB_9_17_port, CI => 
                           SUMB_9_18_port, CO => CARRYB_10_17_port, S => 
                           SUMB_10_17_port);
   S2_10_18 : FA_X1 port map( A => ab_10_18_port, B => CARRYB_9_18_port, CI => 
                           SUMB_9_19_port, CO => CARRYB_10_18_port, S => 
                           SUMB_10_18_port);
   S2_10_19 : FA_X1 port map( A => ab_10_19_port, B => CARRYB_9_19_port, CI => 
                           SUMB_9_20_port, CO => CARRYB_10_19_port, S => 
                           SUMB_10_19_port);
   S2_10_20 : FA_X1 port map( A => ab_10_20_port, B => CARRYB_9_20_port, CI => 
                           SUMB_9_21_port, CO => CARRYB_10_20_port, S => 
                           SUMB_10_20_port);
   S2_10_21 : FA_X1 port map( A => ab_10_21_port, B => CARRYB_9_21_port, CI => 
                           SUMB_9_22_port, CO => n_1054, S => SUMB_10_21_port);
   S1_9_0 : FA_X1 port map( A => ab_9_0_port, B => CARRYB_8_0_port, CI => 
                           SUMB_8_1_port, CO => CARRYB_9_0_port, S => 
                           PRODUCT(9));
   S2_9_1 : FA_X1 port map( A => ab_9_1_port, B => CARRYB_8_1_port, CI => 
                           SUMB_8_2_port, CO => CARRYB_9_1_port, S => 
                           SUMB_9_1_port);
   S2_9_2 : FA_X1 port map( A => ab_9_2_port, B => CARRYB_8_2_port, CI => 
                           SUMB_8_3_port, CO => CARRYB_9_2_port, S => 
                           SUMB_9_2_port);
   S2_9_3 : FA_X1 port map( A => ab_9_3_port, B => CARRYB_8_3_port, CI => 
                           SUMB_8_4_port, CO => CARRYB_9_3_port, S => 
                           SUMB_9_3_port);
   S2_9_4 : FA_X1 port map( A => ab_9_4_port, B => CARRYB_8_4_port, CI => 
                           SUMB_8_5_port, CO => CARRYB_9_4_port, S => 
                           SUMB_9_4_port);
   S2_9_5 : FA_X1 port map( A => ab_9_5_port, B => CARRYB_8_5_port, CI => 
                           SUMB_8_6_port, CO => CARRYB_9_5_port, S => 
                           SUMB_9_5_port);
   S2_9_6 : FA_X1 port map( A => ab_9_6_port, B => CARRYB_8_6_port, CI => 
                           SUMB_8_7_port, CO => CARRYB_9_6_port, S => 
                           SUMB_9_6_port);
   S2_9_7 : FA_X1 port map( A => ab_9_7_port, B => CARRYB_8_7_port, CI => 
                           SUMB_8_8_port, CO => CARRYB_9_7_port, S => 
                           SUMB_9_7_port);
   S2_9_8 : FA_X1 port map( A => ab_9_8_port, B => CARRYB_8_8_port, CI => 
                           SUMB_8_9_port, CO => CARRYB_9_8_port, S => 
                           SUMB_9_8_port);
   S2_9_9 : FA_X1 port map( A => ab_9_9_port, B => CARRYB_8_9_port, CI => 
                           SUMB_8_10_port, CO => CARRYB_9_9_port, S => 
                           SUMB_9_9_port);
   S2_9_10 : FA_X1 port map( A => ab_9_10_port, B => CARRYB_8_10_port, CI => 
                           SUMB_8_11_port, CO => CARRYB_9_10_port, S => 
                           SUMB_9_10_port);
   S2_9_11 : FA_X1 port map( A => ab_9_11_port, B => CARRYB_8_11_port, CI => 
                           SUMB_8_12_port, CO => CARRYB_9_11_port, S => 
                           SUMB_9_11_port);
   S2_9_12 : FA_X1 port map( A => ab_9_12_port, B => CARRYB_8_12_port, CI => 
                           SUMB_8_13_port, CO => CARRYB_9_12_port, S => 
                           SUMB_9_12_port);
   S2_9_13 : FA_X1 port map( A => ab_9_13_port, B => CARRYB_8_13_port, CI => 
                           SUMB_8_14_port, CO => CARRYB_9_13_port, S => 
                           SUMB_9_13_port);
   S2_9_14 : FA_X1 port map( A => ab_9_14_port, B => CARRYB_8_14_port, CI => 
                           SUMB_8_15_port, CO => CARRYB_9_14_port, S => 
                           SUMB_9_14_port);
   S2_9_15 : FA_X1 port map( A => ab_9_15_port, B => CARRYB_8_15_port, CI => 
                           SUMB_8_16_port, CO => CARRYB_9_15_port, S => 
                           SUMB_9_15_port);
   S2_9_16 : FA_X1 port map( A => ab_9_16_port, B => CARRYB_8_16_port, CI => 
                           SUMB_8_17_port, CO => CARRYB_9_16_port, S => 
                           SUMB_9_16_port);
   S2_9_17 : FA_X1 port map( A => ab_9_17_port, B => CARRYB_8_17_port, CI => 
                           SUMB_8_18_port, CO => CARRYB_9_17_port, S => 
                           SUMB_9_17_port);
   S2_9_18 : FA_X1 port map( A => ab_9_18_port, B => CARRYB_8_18_port, CI => 
                           SUMB_8_19_port, CO => CARRYB_9_18_port, S => 
                           SUMB_9_18_port);
   S2_9_19 : FA_X1 port map( A => ab_9_19_port, B => CARRYB_8_19_port, CI => 
                           SUMB_8_20_port, CO => CARRYB_9_19_port, S => 
                           SUMB_9_19_port);
   S2_9_20 : FA_X1 port map( A => ab_9_20_port, B => CARRYB_8_20_port, CI => 
                           SUMB_8_21_port, CO => CARRYB_9_20_port, S => 
                           SUMB_9_20_port);
   S2_9_21 : FA_X1 port map( A => ab_9_21_port, B => CARRYB_8_21_port, CI => 
                           SUMB_8_22_port, CO => CARRYB_9_21_port, S => 
                           SUMB_9_21_port);
   S2_9_22 : FA_X1 port map( A => ab_9_22_port, B => CARRYB_8_22_port, CI => 
                           SUMB_8_23_port, CO => n_1055, S => SUMB_9_22_port);
   S1_8_0 : FA_X1 port map( A => ab_8_0_port, B => CARRYB_7_0_port, CI => 
                           SUMB_7_1_port, CO => CARRYB_8_0_port, S => 
                           PRODUCT(8));
   S2_8_1 : FA_X1 port map( A => ab_8_1_port, B => CARRYB_7_1_port, CI => 
                           SUMB_7_2_port, CO => CARRYB_8_1_port, S => 
                           SUMB_8_1_port);
   S2_8_2 : FA_X1 port map( A => ab_8_2_port, B => CARRYB_7_2_port, CI => 
                           SUMB_7_3_port, CO => CARRYB_8_2_port, S => 
                           SUMB_8_2_port);
   S2_8_3 : FA_X1 port map( A => ab_8_3_port, B => CARRYB_7_3_port, CI => 
                           SUMB_7_4_port, CO => CARRYB_8_3_port, S => 
                           SUMB_8_3_port);
   S2_8_4 : FA_X1 port map( A => ab_8_4_port, B => CARRYB_7_4_port, CI => 
                           SUMB_7_5_port, CO => CARRYB_8_4_port, S => 
                           SUMB_8_4_port);
   S2_8_5 : FA_X1 port map( A => ab_8_5_port, B => CARRYB_7_5_port, CI => 
                           SUMB_7_6_port, CO => CARRYB_8_5_port, S => 
                           SUMB_8_5_port);
   S2_8_6 : FA_X1 port map( A => ab_8_6_port, B => CARRYB_7_6_port, CI => 
                           SUMB_7_7_port, CO => CARRYB_8_6_port, S => 
                           SUMB_8_6_port);
   S2_8_7 : FA_X1 port map( A => ab_8_7_port, B => CARRYB_7_7_port, CI => 
                           SUMB_7_8_port, CO => CARRYB_8_7_port, S => 
                           SUMB_8_7_port);
   S2_8_8 : FA_X1 port map( A => ab_8_8_port, B => CARRYB_7_8_port, CI => 
                           SUMB_7_9_port, CO => CARRYB_8_8_port, S => 
                           SUMB_8_8_port);
   S2_8_9 : FA_X1 port map( A => ab_8_9_port, B => CARRYB_7_9_port, CI => 
                           SUMB_7_10_port, CO => CARRYB_8_9_port, S => 
                           SUMB_8_9_port);
   S2_8_10 : FA_X1 port map( A => ab_8_10_port, B => CARRYB_7_10_port, CI => 
                           SUMB_7_11_port, CO => CARRYB_8_10_port, S => 
                           SUMB_8_10_port);
   S2_8_11 : FA_X1 port map( A => ab_8_11_port, B => CARRYB_7_11_port, CI => 
                           SUMB_7_12_port, CO => CARRYB_8_11_port, S => 
                           SUMB_8_11_port);
   S2_8_12 : FA_X1 port map( A => ab_8_12_port, B => CARRYB_7_12_port, CI => 
                           SUMB_7_13_port, CO => CARRYB_8_12_port, S => 
                           SUMB_8_12_port);
   S2_8_13 : FA_X1 port map( A => ab_8_13_port, B => CARRYB_7_13_port, CI => 
                           SUMB_7_14_port, CO => CARRYB_8_13_port, S => 
                           SUMB_8_13_port);
   S2_8_14 : FA_X1 port map( A => ab_8_14_port, B => CARRYB_7_14_port, CI => 
                           SUMB_7_15_port, CO => CARRYB_8_14_port, S => 
                           SUMB_8_14_port);
   S2_8_15 : FA_X1 port map( A => ab_8_15_port, B => CARRYB_7_15_port, CI => 
                           SUMB_7_16_port, CO => CARRYB_8_15_port, S => 
                           SUMB_8_15_port);
   S2_8_16 : FA_X1 port map( A => ab_8_16_port, B => CARRYB_7_16_port, CI => 
                           SUMB_7_17_port, CO => CARRYB_8_16_port, S => 
                           SUMB_8_16_port);
   S2_8_17 : FA_X1 port map( A => ab_8_17_port, B => CARRYB_7_17_port, CI => 
                           SUMB_7_18_port, CO => CARRYB_8_17_port, S => 
                           SUMB_8_17_port);
   S2_8_18 : FA_X1 port map( A => ab_8_18_port, B => CARRYB_7_18_port, CI => 
                           SUMB_7_19_port, CO => CARRYB_8_18_port, S => 
                           SUMB_8_18_port);
   S2_8_19 : FA_X1 port map( A => ab_8_19_port, B => CARRYB_7_19_port, CI => 
                           SUMB_7_20_port, CO => CARRYB_8_19_port, S => 
                           SUMB_8_19_port);
   S2_8_20 : FA_X1 port map( A => ab_8_20_port, B => CARRYB_7_20_port, CI => 
                           SUMB_7_21_port, CO => CARRYB_8_20_port, S => 
                           SUMB_8_20_port);
   S2_8_21 : FA_X1 port map( A => ab_8_21_port, B => CARRYB_7_21_port, CI => 
                           SUMB_7_22_port, CO => CARRYB_8_21_port, S => 
                           SUMB_8_21_port);
   S2_8_22 : FA_X1 port map( A => ab_8_22_port, B => CARRYB_7_22_port, CI => 
                           SUMB_7_23_port, CO => CARRYB_8_22_port, S => 
                           SUMB_8_22_port);
   S2_8_23 : FA_X1 port map( A => ab_8_23_port, B => CARRYB_7_23_port, CI => 
                           SUMB_7_24_port, CO => n_1056, S => SUMB_8_23_port);
   S1_7_0 : FA_X1 port map( A => ab_7_0_port, B => CARRYB_6_0_port, CI => 
                           SUMB_6_1_port, CO => CARRYB_7_0_port, S => 
                           PRODUCT(7));
   S2_7_1 : FA_X1 port map( A => ab_7_1_port, B => CARRYB_6_1_port, CI => 
                           SUMB_6_2_port, CO => CARRYB_7_1_port, S => 
                           SUMB_7_1_port);
   S2_7_2 : FA_X1 port map( A => ab_7_2_port, B => CARRYB_6_2_port, CI => 
                           SUMB_6_3_port, CO => CARRYB_7_2_port, S => 
                           SUMB_7_2_port);
   S2_7_3 : FA_X1 port map( A => ab_7_3_port, B => CARRYB_6_3_port, CI => 
                           SUMB_6_4_port, CO => CARRYB_7_3_port, S => 
                           SUMB_7_3_port);
   S2_7_4 : FA_X1 port map( A => ab_7_4_port, B => CARRYB_6_4_port, CI => 
                           SUMB_6_5_port, CO => CARRYB_7_4_port, S => 
                           SUMB_7_4_port);
   S2_7_5 : FA_X1 port map( A => ab_7_5_port, B => CARRYB_6_5_port, CI => 
                           SUMB_6_6_port, CO => CARRYB_7_5_port, S => 
                           SUMB_7_5_port);
   S2_7_6 : FA_X1 port map( A => ab_7_6_port, B => CARRYB_6_6_port, CI => 
                           SUMB_6_7_port, CO => CARRYB_7_6_port, S => 
                           SUMB_7_6_port);
   S2_7_7 : FA_X1 port map( A => ab_7_7_port, B => CARRYB_6_7_port, CI => 
                           SUMB_6_8_port, CO => CARRYB_7_7_port, S => 
                           SUMB_7_7_port);
   S2_7_8 : FA_X1 port map( A => ab_7_8_port, B => CARRYB_6_8_port, CI => 
                           SUMB_6_9_port, CO => CARRYB_7_8_port, S => 
                           SUMB_7_8_port);
   S2_7_9 : FA_X1 port map( A => ab_7_9_port, B => CARRYB_6_9_port, CI => 
                           SUMB_6_10_port, CO => CARRYB_7_9_port, S => 
                           SUMB_7_9_port);
   S2_7_10 : FA_X1 port map( A => ab_7_10_port, B => CARRYB_6_10_port, CI => 
                           SUMB_6_11_port, CO => CARRYB_7_10_port, S => 
                           SUMB_7_10_port);
   S2_7_11 : FA_X1 port map( A => ab_7_11_port, B => CARRYB_6_11_port, CI => 
                           SUMB_6_12_port, CO => CARRYB_7_11_port, S => 
                           SUMB_7_11_port);
   S2_7_12 : FA_X1 port map( A => ab_7_12_port, B => CARRYB_6_12_port, CI => 
                           SUMB_6_13_port, CO => CARRYB_7_12_port, S => 
                           SUMB_7_12_port);
   S2_7_13 : FA_X1 port map( A => ab_7_13_port, B => CARRYB_6_13_port, CI => 
                           SUMB_6_14_port, CO => CARRYB_7_13_port, S => 
                           SUMB_7_13_port);
   S2_7_14 : FA_X1 port map( A => ab_7_14_port, B => CARRYB_6_14_port, CI => 
                           SUMB_6_15_port, CO => CARRYB_7_14_port, S => 
                           SUMB_7_14_port);
   S2_7_15 : FA_X1 port map( A => ab_7_15_port, B => CARRYB_6_15_port, CI => 
                           SUMB_6_16_port, CO => CARRYB_7_15_port, S => 
                           SUMB_7_15_port);
   S2_7_16 : FA_X1 port map( A => ab_7_16_port, B => CARRYB_6_16_port, CI => 
                           SUMB_6_17_port, CO => CARRYB_7_16_port, S => 
                           SUMB_7_16_port);
   S2_7_17 : FA_X1 port map( A => ab_7_17_port, B => CARRYB_6_17_port, CI => 
                           SUMB_6_18_port, CO => CARRYB_7_17_port, S => 
                           SUMB_7_17_port);
   S2_7_18 : FA_X1 port map( A => ab_7_18_port, B => CARRYB_6_18_port, CI => 
                           SUMB_6_19_port, CO => CARRYB_7_18_port, S => 
                           SUMB_7_18_port);
   S2_7_19 : FA_X1 port map( A => ab_7_19_port, B => CARRYB_6_19_port, CI => 
                           SUMB_6_20_port, CO => CARRYB_7_19_port, S => 
                           SUMB_7_19_port);
   S2_7_20 : FA_X1 port map( A => ab_7_20_port, B => CARRYB_6_20_port, CI => 
                           SUMB_6_21_port, CO => CARRYB_7_20_port, S => 
                           SUMB_7_20_port);
   S2_7_21 : FA_X1 port map( A => ab_7_21_port, B => CARRYB_6_21_port, CI => 
                           SUMB_6_22_port, CO => CARRYB_7_21_port, S => 
                           SUMB_7_21_port);
   S2_7_22 : FA_X1 port map( A => ab_7_22_port, B => CARRYB_6_22_port, CI => 
                           SUMB_6_23_port, CO => CARRYB_7_22_port, S => 
                           SUMB_7_22_port);
   S2_7_23 : FA_X1 port map( A => ab_7_23_port, B => CARRYB_6_23_port, CI => 
                           SUMB_6_24_port, CO => CARRYB_7_23_port, S => 
                           SUMB_7_23_port);
   S2_7_24 : FA_X1 port map( A => ab_7_24_port, B => CARRYB_6_24_port, CI => 
                           SUMB_6_25_port, CO => n_1057, S => SUMB_7_24_port);
   S1_6_0 : FA_X1 port map( A => ab_6_0_port, B => CARRYB_5_0_port, CI => 
                           SUMB_5_1_port, CO => CARRYB_6_0_port, S => 
                           PRODUCT(6));
   S2_6_1 : FA_X1 port map( A => ab_6_1_port, B => CARRYB_5_1_port, CI => 
                           SUMB_5_2_port, CO => CARRYB_6_1_port, S => 
                           SUMB_6_1_port);
   S2_6_2 : FA_X1 port map( A => ab_6_2_port, B => CARRYB_5_2_port, CI => 
                           SUMB_5_3_port, CO => CARRYB_6_2_port, S => 
                           SUMB_6_2_port);
   S2_6_3 : FA_X1 port map( A => ab_6_3_port, B => CARRYB_5_3_port, CI => 
                           SUMB_5_4_port, CO => CARRYB_6_3_port, S => 
                           SUMB_6_3_port);
   S2_6_4 : FA_X1 port map( A => ab_6_4_port, B => CARRYB_5_4_port, CI => 
                           SUMB_5_5_port, CO => CARRYB_6_4_port, S => 
                           SUMB_6_4_port);
   S2_6_5 : FA_X1 port map( A => ab_6_5_port, B => CARRYB_5_5_port, CI => 
                           SUMB_5_6_port, CO => CARRYB_6_5_port, S => 
                           SUMB_6_5_port);
   S2_6_6 : FA_X1 port map( A => ab_6_6_port, B => CARRYB_5_6_port, CI => 
                           SUMB_5_7_port, CO => CARRYB_6_6_port, S => 
                           SUMB_6_6_port);
   S2_6_7 : FA_X1 port map( A => ab_6_7_port, B => CARRYB_5_7_port, CI => 
                           SUMB_5_8_port, CO => CARRYB_6_7_port, S => 
                           SUMB_6_7_port);
   S2_6_8 : FA_X1 port map( A => ab_6_8_port, B => CARRYB_5_8_port, CI => 
                           SUMB_5_9_port, CO => CARRYB_6_8_port, S => 
                           SUMB_6_8_port);
   S2_6_9 : FA_X1 port map( A => ab_6_9_port, B => CARRYB_5_9_port, CI => 
                           SUMB_5_10_port, CO => CARRYB_6_9_port, S => 
                           SUMB_6_9_port);
   S2_6_10 : FA_X1 port map( A => ab_6_10_port, B => CARRYB_5_10_port, CI => 
                           SUMB_5_11_port, CO => CARRYB_6_10_port, S => 
                           SUMB_6_10_port);
   S2_6_11 : FA_X1 port map( A => ab_6_11_port, B => CARRYB_5_11_port, CI => 
                           SUMB_5_12_port, CO => CARRYB_6_11_port, S => 
                           SUMB_6_11_port);
   S2_6_12 : FA_X1 port map( A => ab_6_12_port, B => CARRYB_5_12_port, CI => 
                           SUMB_5_13_port, CO => CARRYB_6_12_port, S => 
                           SUMB_6_12_port);
   S2_6_13 : FA_X1 port map( A => ab_6_13_port, B => CARRYB_5_13_port, CI => 
                           SUMB_5_14_port, CO => CARRYB_6_13_port, S => 
                           SUMB_6_13_port);
   S2_6_14 : FA_X1 port map( A => ab_6_14_port, B => CARRYB_5_14_port, CI => 
                           SUMB_5_15_port, CO => CARRYB_6_14_port, S => 
                           SUMB_6_14_port);
   S2_6_15 : FA_X1 port map( A => ab_6_15_port, B => CARRYB_5_15_port, CI => 
                           SUMB_5_16_port, CO => CARRYB_6_15_port, S => 
                           SUMB_6_15_port);
   S2_6_16 : FA_X1 port map( A => ab_6_16_port, B => CARRYB_5_16_port, CI => 
                           SUMB_5_17_port, CO => CARRYB_6_16_port, S => 
                           SUMB_6_16_port);
   S2_6_17 : FA_X1 port map( A => ab_6_17_port, B => CARRYB_5_17_port, CI => 
                           SUMB_5_18_port, CO => CARRYB_6_17_port, S => 
                           SUMB_6_17_port);
   S2_6_18 : FA_X1 port map( A => ab_6_18_port, B => CARRYB_5_18_port, CI => 
                           SUMB_5_19_port, CO => CARRYB_6_18_port, S => 
                           SUMB_6_18_port);
   S2_6_19 : FA_X1 port map( A => ab_6_19_port, B => CARRYB_5_19_port, CI => 
                           SUMB_5_20_port, CO => CARRYB_6_19_port, S => 
                           SUMB_6_19_port);
   S2_6_20 : FA_X1 port map( A => ab_6_20_port, B => CARRYB_5_20_port, CI => 
                           SUMB_5_21_port, CO => CARRYB_6_20_port, S => 
                           SUMB_6_20_port);
   S2_6_21 : FA_X1 port map( A => ab_6_21_port, B => CARRYB_5_21_port, CI => 
                           SUMB_5_22_port, CO => CARRYB_6_21_port, S => 
                           SUMB_6_21_port);
   S2_6_22 : FA_X1 port map( A => ab_6_22_port, B => CARRYB_5_22_port, CI => 
                           SUMB_5_23_port, CO => CARRYB_6_22_port, S => 
                           SUMB_6_22_port);
   S2_6_23 : FA_X1 port map( A => ab_6_23_port, B => CARRYB_5_23_port, CI => 
                           SUMB_5_24_port, CO => CARRYB_6_23_port, S => 
                           SUMB_6_23_port);
   S2_6_24 : FA_X1 port map( A => ab_6_24_port, B => CARRYB_5_24_port, CI => 
                           SUMB_5_25_port, CO => CARRYB_6_24_port, S => 
                           SUMB_6_24_port);
   S2_6_25 : FA_X1 port map( A => ab_6_25_port, B => CARRYB_5_25_port, CI => 
                           SUMB_5_26_port, CO => n_1058, S => SUMB_6_25_port);
   S1_5_0 : FA_X1 port map( A => ab_5_0_port, B => CARRYB_4_0_port, CI => 
                           SUMB_4_1_port, CO => CARRYB_5_0_port, S => 
                           PRODUCT(5));
   S2_5_1 : FA_X1 port map( A => ab_5_1_port, B => CARRYB_4_1_port, CI => 
                           SUMB_4_2_port, CO => CARRYB_5_1_port, S => 
                           SUMB_5_1_port);
   S2_5_2 : FA_X1 port map( A => ab_5_2_port, B => CARRYB_4_2_port, CI => 
                           SUMB_4_3_port, CO => CARRYB_5_2_port, S => 
                           SUMB_5_2_port);
   S2_5_3 : FA_X1 port map( A => ab_5_3_port, B => CARRYB_4_3_port, CI => 
                           SUMB_4_4_port, CO => CARRYB_5_3_port, S => 
                           SUMB_5_3_port);
   S2_5_4 : FA_X1 port map( A => ab_5_4_port, B => CARRYB_4_4_port, CI => 
                           SUMB_4_5_port, CO => CARRYB_5_4_port, S => 
                           SUMB_5_4_port);
   S2_5_5 : FA_X1 port map( A => ab_5_5_port, B => CARRYB_4_5_port, CI => 
                           SUMB_4_6_port, CO => CARRYB_5_5_port, S => 
                           SUMB_5_5_port);
   S2_5_6 : FA_X1 port map( A => ab_5_6_port, B => CARRYB_4_6_port, CI => 
                           SUMB_4_7_port, CO => CARRYB_5_6_port, S => 
                           SUMB_5_6_port);
   S2_5_7 : FA_X1 port map( A => ab_5_7_port, B => CARRYB_4_7_port, CI => 
                           SUMB_4_8_port, CO => CARRYB_5_7_port, S => 
                           SUMB_5_7_port);
   S2_5_8 : FA_X1 port map( A => ab_5_8_port, B => CARRYB_4_8_port, CI => 
                           SUMB_4_9_port, CO => CARRYB_5_8_port, S => 
                           SUMB_5_8_port);
   S2_5_9 : FA_X1 port map( A => ab_5_9_port, B => CARRYB_4_9_port, CI => 
                           SUMB_4_10_port, CO => CARRYB_5_9_port, S => 
                           SUMB_5_9_port);
   S2_5_10 : FA_X1 port map( A => ab_5_10_port, B => CARRYB_4_10_port, CI => 
                           SUMB_4_11_port, CO => CARRYB_5_10_port, S => 
                           SUMB_5_10_port);
   S2_5_11 : FA_X1 port map( A => ab_5_11_port, B => CARRYB_4_11_port, CI => 
                           SUMB_4_12_port, CO => CARRYB_5_11_port, S => 
                           SUMB_5_11_port);
   S2_5_12 : FA_X1 port map( A => ab_5_12_port, B => CARRYB_4_12_port, CI => 
                           SUMB_4_13_port, CO => CARRYB_5_12_port, S => 
                           SUMB_5_12_port);
   S2_5_13 : FA_X1 port map( A => ab_5_13_port, B => CARRYB_4_13_port, CI => 
                           SUMB_4_14_port, CO => CARRYB_5_13_port, S => 
                           SUMB_5_13_port);
   S2_5_14 : FA_X1 port map( A => ab_5_14_port, B => CARRYB_4_14_port, CI => 
                           SUMB_4_15_port, CO => CARRYB_5_14_port, S => 
                           SUMB_5_14_port);
   S2_5_15 : FA_X1 port map( A => ab_5_15_port, B => CARRYB_4_15_port, CI => 
                           SUMB_4_16_port, CO => CARRYB_5_15_port, S => 
                           SUMB_5_15_port);
   S2_5_16 : FA_X1 port map( A => ab_5_16_port, B => CARRYB_4_16_port, CI => 
                           SUMB_4_17_port, CO => CARRYB_5_16_port, S => 
                           SUMB_5_16_port);
   S2_5_17 : FA_X1 port map( A => ab_5_17_port, B => CARRYB_4_17_port, CI => 
                           SUMB_4_18_port, CO => CARRYB_5_17_port, S => 
                           SUMB_5_17_port);
   S2_5_18 : FA_X1 port map( A => ab_5_18_port, B => CARRYB_4_18_port, CI => 
                           SUMB_4_19_port, CO => CARRYB_5_18_port, S => 
                           SUMB_5_18_port);
   S2_5_19 : FA_X1 port map( A => ab_5_19_port, B => CARRYB_4_19_port, CI => 
                           SUMB_4_20_port, CO => CARRYB_5_19_port, S => 
                           SUMB_5_19_port);
   S2_5_20 : FA_X1 port map( A => ab_5_20_port, B => CARRYB_4_20_port, CI => 
                           SUMB_4_21_port, CO => CARRYB_5_20_port, S => 
                           SUMB_5_20_port);
   S2_5_21 : FA_X1 port map( A => ab_5_21_port, B => CARRYB_4_21_port, CI => 
                           SUMB_4_22_port, CO => CARRYB_5_21_port, S => 
                           SUMB_5_21_port);
   S2_5_22 : FA_X1 port map( A => ab_5_22_port, B => CARRYB_4_22_port, CI => 
                           SUMB_4_23_port, CO => CARRYB_5_22_port, S => 
                           SUMB_5_22_port);
   S2_5_23 : FA_X1 port map( A => ab_5_23_port, B => CARRYB_4_23_port, CI => 
                           SUMB_4_24_port, CO => CARRYB_5_23_port, S => 
                           SUMB_5_23_port);
   S2_5_24 : FA_X1 port map( A => ab_5_24_port, B => CARRYB_4_24_port, CI => 
                           SUMB_4_25_port, CO => CARRYB_5_24_port, S => 
                           SUMB_5_24_port);
   S2_5_25 : FA_X1 port map( A => ab_5_25_port, B => CARRYB_4_25_port, CI => 
                           SUMB_4_26_port, CO => CARRYB_5_25_port, S => 
                           SUMB_5_25_port);
   S2_5_26 : FA_X1 port map( A => ab_5_26_port, B => CARRYB_4_26_port, CI => 
                           SUMB_4_27_port, CO => n_1059, S => SUMB_5_26_port);
   S1_4_0 : FA_X1 port map( A => ab_4_0_port, B => CARRYB_3_0_port, CI => 
                           SUMB_3_1_port, CO => CARRYB_4_0_port, S => 
                           PRODUCT(4));
   S2_4_1 : FA_X1 port map( A => ab_4_1_port, B => CARRYB_3_1_port, CI => 
                           SUMB_3_2_port, CO => CARRYB_4_1_port, S => 
                           SUMB_4_1_port);
   S2_4_2 : FA_X1 port map( A => ab_4_2_port, B => CARRYB_3_2_port, CI => 
                           SUMB_3_3_port, CO => CARRYB_4_2_port, S => 
                           SUMB_4_2_port);
   S2_4_3 : FA_X1 port map( A => ab_4_3_port, B => CARRYB_3_3_port, CI => 
                           SUMB_3_4_port, CO => CARRYB_4_3_port, S => 
                           SUMB_4_3_port);
   S2_4_4 : FA_X1 port map( A => ab_4_4_port, B => CARRYB_3_4_port, CI => 
                           SUMB_3_5_port, CO => CARRYB_4_4_port, S => 
                           SUMB_4_4_port);
   S2_4_5 : FA_X1 port map( A => ab_4_5_port, B => CARRYB_3_5_port, CI => 
                           SUMB_3_6_port, CO => CARRYB_4_5_port, S => 
                           SUMB_4_5_port);
   S2_4_6 : FA_X1 port map( A => ab_4_6_port, B => CARRYB_3_6_port, CI => 
                           SUMB_3_7_port, CO => CARRYB_4_6_port, S => 
                           SUMB_4_6_port);
   S2_4_7 : FA_X1 port map( A => ab_4_7_port, B => CARRYB_3_7_port, CI => 
                           SUMB_3_8_port, CO => CARRYB_4_7_port, S => 
                           SUMB_4_7_port);
   S2_4_8 : FA_X1 port map( A => ab_4_8_port, B => CARRYB_3_8_port, CI => 
                           SUMB_3_9_port, CO => CARRYB_4_8_port, S => 
                           SUMB_4_8_port);
   S2_4_9 : FA_X1 port map( A => ab_4_9_port, B => CARRYB_3_9_port, CI => 
                           SUMB_3_10_port, CO => CARRYB_4_9_port, S => 
                           SUMB_4_9_port);
   S2_4_10 : FA_X1 port map( A => ab_4_10_port, B => CARRYB_3_10_port, CI => 
                           SUMB_3_11_port, CO => CARRYB_4_10_port, S => 
                           SUMB_4_10_port);
   S2_4_11 : FA_X1 port map( A => ab_4_11_port, B => CARRYB_3_11_port, CI => 
                           SUMB_3_12_port, CO => CARRYB_4_11_port, S => 
                           SUMB_4_11_port);
   S2_4_12 : FA_X1 port map( A => ab_4_12_port, B => CARRYB_3_12_port, CI => 
                           SUMB_3_13_port, CO => CARRYB_4_12_port, S => 
                           SUMB_4_12_port);
   S2_4_13 : FA_X1 port map( A => ab_4_13_port, B => CARRYB_3_13_port, CI => 
                           SUMB_3_14_port, CO => CARRYB_4_13_port, S => 
                           SUMB_4_13_port);
   S2_4_14 : FA_X1 port map( A => ab_4_14_port, B => CARRYB_3_14_port, CI => 
                           SUMB_3_15_port, CO => CARRYB_4_14_port, S => 
                           SUMB_4_14_port);
   S2_4_15 : FA_X1 port map( A => ab_4_15_port, B => CARRYB_3_15_port, CI => 
                           SUMB_3_16_port, CO => CARRYB_4_15_port, S => 
                           SUMB_4_15_port);
   S2_4_16 : FA_X1 port map( A => ab_4_16_port, B => CARRYB_3_16_port, CI => 
                           SUMB_3_17_port, CO => CARRYB_4_16_port, S => 
                           SUMB_4_16_port);
   S2_4_17 : FA_X1 port map( A => ab_4_17_port, B => CARRYB_3_17_port, CI => 
                           SUMB_3_18_port, CO => CARRYB_4_17_port, S => 
                           SUMB_4_17_port);
   S2_4_18 : FA_X1 port map( A => ab_4_18_port, B => CARRYB_3_18_port, CI => 
                           SUMB_3_19_port, CO => CARRYB_4_18_port, S => 
                           SUMB_4_18_port);
   S2_4_19 : FA_X1 port map( A => ab_4_19_port, B => CARRYB_3_19_port, CI => 
                           SUMB_3_20_port, CO => CARRYB_4_19_port, S => 
                           SUMB_4_19_port);
   S2_4_20 : FA_X1 port map( A => ab_4_20_port, B => CARRYB_3_20_port, CI => 
                           SUMB_3_21_port, CO => CARRYB_4_20_port, S => 
                           SUMB_4_20_port);
   S2_4_21 : FA_X1 port map( A => ab_4_21_port, B => CARRYB_3_21_port, CI => 
                           SUMB_3_22_port, CO => CARRYB_4_21_port, S => 
                           SUMB_4_21_port);
   S2_4_22 : FA_X1 port map( A => ab_4_22_port, B => CARRYB_3_22_port, CI => 
                           SUMB_3_23_port, CO => CARRYB_4_22_port, S => 
                           SUMB_4_22_port);
   S2_4_23 : FA_X1 port map( A => ab_4_23_port, B => CARRYB_3_23_port, CI => 
                           SUMB_3_24_port, CO => CARRYB_4_23_port, S => 
                           SUMB_4_23_port);
   S2_4_24 : FA_X1 port map( A => ab_4_24_port, B => CARRYB_3_24_port, CI => 
                           SUMB_3_25_port, CO => CARRYB_4_24_port, S => 
                           SUMB_4_24_port);
   S2_4_25 : FA_X1 port map( A => ab_4_25_port, B => CARRYB_3_25_port, CI => 
                           SUMB_3_26_port, CO => CARRYB_4_25_port, S => 
                           SUMB_4_25_port);
   S2_4_26 : FA_X1 port map( A => ab_4_26_port, B => CARRYB_3_26_port, CI => 
                           SUMB_3_27_port, CO => CARRYB_4_26_port, S => 
                           SUMB_4_26_port);
   S2_4_27 : FA_X1 port map( A => ab_4_27_port, B => CARRYB_3_27_port, CI => 
                           SUMB_3_28_port, CO => n_1060, S => SUMB_4_27_port);
   S1_3_0 : FA_X1 port map( A => ab_3_0_port, B => CARRYB_2_0_port, CI => 
                           SUMB_2_1_port, CO => CARRYB_3_0_port, S => 
                           PRODUCT(3));
   S2_3_1 : FA_X1 port map( A => ab_3_1_port, B => CARRYB_2_1_port, CI => 
                           SUMB_2_2_port, CO => CARRYB_3_1_port, S => 
                           SUMB_3_1_port);
   S2_3_2 : FA_X1 port map( A => ab_3_2_port, B => CARRYB_2_2_port, CI => 
                           SUMB_2_3_port, CO => CARRYB_3_2_port, S => 
                           SUMB_3_2_port);
   S2_3_3 : FA_X1 port map( A => ab_3_3_port, B => CARRYB_2_3_port, CI => 
                           SUMB_2_4_port, CO => CARRYB_3_3_port, S => 
                           SUMB_3_3_port);
   S2_3_4 : FA_X1 port map( A => ab_3_4_port, B => CARRYB_2_4_port, CI => 
                           SUMB_2_5_port, CO => CARRYB_3_4_port, S => 
                           SUMB_3_4_port);
   S2_3_5 : FA_X1 port map( A => ab_3_5_port, B => CARRYB_2_5_port, CI => 
                           SUMB_2_6_port, CO => CARRYB_3_5_port, S => 
                           SUMB_3_5_port);
   S2_3_6 : FA_X1 port map( A => ab_3_6_port, B => CARRYB_2_6_port, CI => 
                           SUMB_2_7_port, CO => CARRYB_3_6_port, S => 
                           SUMB_3_6_port);
   S2_3_7 : FA_X1 port map( A => ab_3_7_port, B => CARRYB_2_7_port, CI => 
                           SUMB_2_8_port, CO => CARRYB_3_7_port, S => 
                           SUMB_3_7_port);
   S2_3_8 : FA_X1 port map( A => ab_3_8_port, B => CARRYB_2_8_port, CI => 
                           SUMB_2_9_port, CO => CARRYB_3_8_port, S => 
                           SUMB_3_8_port);
   S2_3_9 : FA_X1 port map( A => ab_3_9_port, B => CARRYB_2_9_port, CI => 
                           SUMB_2_10_port, CO => CARRYB_3_9_port, S => 
                           SUMB_3_9_port);
   S2_3_10 : FA_X1 port map( A => ab_3_10_port, B => CARRYB_2_10_port, CI => 
                           SUMB_2_11_port, CO => CARRYB_3_10_port, S => 
                           SUMB_3_10_port);
   S2_3_11 : FA_X1 port map( A => ab_3_11_port, B => CARRYB_2_11_port, CI => 
                           SUMB_2_12_port, CO => CARRYB_3_11_port, S => 
                           SUMB_3_11_port);
   S2_3_12 : FA_X1 port map( A => ab_3_12_port, B => CARRYB_2_12_port, CI => 
                           SUMB_2_13_port, CO => CARRYB_3_12_port, S => 
                           SUMB_3_12_port);
   S2_3_13 : FA_X1 port map( A => ab_3_13_port, B => CARRYB_2_13_port, CI => 
                           SUMB_2_14_port, CO => CARRYB_3_13_port, S => 
                           SUMB_3_13_port);
   S2_3_14 : FA_X1 port map( A => ab_3_14_port, B => CARRYB_2_14_port, CI => 
                           SUMB_2_15_port, CO => CARRYB_3_14_port, S => 
                           SUMB_3_14_port);
   S2_3_15 : FA_X1 port map( A => ab_3_15_port, B => CARRYB_2_15_port, CI => 
                           SUMB_2_16_port, CO => CARRYB_3_15_port, S => 
                           SUMB_3_15_port);
   S2_3_16 : FA_X1 port map( A => ab_3_16_port, B => CARRYB_2_16_port, CI => 
                           SUMB_2_17_port, CO => CARRYB_3_16_port, S => 
                           SUMB_3_16_port);
   S2_3_17 : FA_X1 port map( A => ab_3_17_port, B => CARRYB_2_17_port, CI => 
                           SUMB_2_18_port, CO => CARRYB_3_17_port, S => 
                           SUMB_3_17_port);
   S2_3_18 : FA_X1 port map( A => ab_3_18_port, B => CARRYB_2_18_port, CI => 
                           SUMB_2_19_port, CO => CARRYB_3_18_port, S => 
                           SUMB_3_18_port);
   S2_3_19 : FA_X1 port map( A => ab_3_19_port, B => CARRYB_2_19_port, CI => 
                           SUMB_2_20_port, CO => CARRYB_3_19_port, S => 
                           SUMB_3_19_port);
   S2_3_20 : FA_X1 port map( A => ab_3_20_port, B => CARRYB_2_20_port, CI => 
                           SUMB_2_21_port, CO => CARRYB_3_20_port, S => 
                           SUMB_3_20_port);
   S2_3_21 : FA_X1 port map( A => ab_3_21_port, B => CARRYB_2_21_port, CI => 
                           SUMB_2_22_port, CO => CARRYB_3_21_port, S => 
                           SUMB_3_21_port);
   S2_3_22 : FA_X1 port map( A => ab_3_22_port, B => CARRYB_2_22_port, CI => 
                           SUMB_2_23_port, CO => CARRYB_3_22_port, S => 
                           SUMB_3_22_port);
   S2_3_23 : FA_X1 port map( A => ab_3_23_port, B => CARRYB_2_23_port, CI => 
                           SUMB_2_24_port, CO => CARRYB_3_23_port, S => 
                           SUMB_3_23_port);
   S2_3_24 : FA_X1 port map( A => ab_3_24_port, B => CARRYB_2_24_port, CI => 
                           SUMB_2_25_port, CO => CARRYB_3_24_port, S => 
                           SUMB_3_24_port);
   S2_3_25 : FA_X1 port map( A => ab_3_25_port, B => CARRYB_2_25_port, CI => 
                           SUMB_2_26_port, CO => CARRYB_3_25_port, S => 
                           SUMB_3_25_port);
   S2_3_26 : FA_X1 port map( A => ab_3_26_port, B => CARRYB_2_26_port, CI => 
                           SUMB_2_27_port, CO => CARRYB_3_26_port, S => 
                           SUMB_3_26_port);
   S2_3_27 : FA_X1 port map( A => ab_3_27_port, B => CARRYB_2_27_port, CI => 
                           SUMB_2_28_port, CO => CARRYB_3_27_port, S => 
                           SUMB_3_27_port);
   S2_3_28 : FA_X1 port map( A => ab_3_28_port, B => CARRYB_2_28_port, CI => 
                           SUMB_2_29_port, CO => n_1061, S => SUMB_3_28_port);
   S1_2_0 : FA_X1 port map( A => ab_2_0_port, B => n24, CI => n53, CO => 
                           CARRYB_2_0_port, S => PRODUCT(2));
   S2_2_1 : FA_X1 port map( A => ab_2_1_port, B => n23, CI => n59, CO => 
                           CARRYB_2_1_port, S => SUMB_2_1_port);
   S2_2_2 : FA_X1 port map( A => ab_2_2_port, B => n30, CI => n58, CO => 
                           CARRYB_2_2_port, S => SUMB_2_2_port);
   S2_2_3 : FA_X1 port map( A => ab_2_3_port, B => n29, CI => n57, CO => 
                           CARRYB_2_3_port, S => SUMB_2_3_port);
   S2_2_4 : FA_X1 port map( A => ab_2_4_port, B => n28, CI => n56, CO => 
                           CARRYB_2_4_port, S => SUMB_2_4_port);
   S2_2_5 : FA_X1 port map( A => ab_2_5_port, B => n27, CI => n55, CO => 
                           CARRYB_2_5_port, S => SUMB_2_5_port);
   S2_2_6 : FA_X1 port map( A => ab_2_6_port, B => n26, CI => n54, CO => 
                           CARRYB_2_6_port, S => SUMB_2_6_port);
   S2_2_7 : FA_X1 port map( A => ab_2_7_port, B => n25, CI => n50, CO => 
                           CARRYB_2_7_port, S => SUMB_2_7_port);
   S2_2_8 : FA_X1 port map( A => ab_2_8_port, B => n21, CI => n51, CO => 
                           CARRYB_2_8_port, S => SUMB_2_8_port);
   S2_2_9 : FA_X1 port map( A => ab_2_9_port, B => n22, CI => n52, CO => 
                           CARRYB_2_9_port, S => SUMB_2_9_port);
   S2_2_10 : FA_X1 port map( A => ab_2_10_port, B => n49, CI => n20, CO => 
                           CARRYB_2_10_port, S => SUMB_2_10_port);
   S2_2_11 : FA_X1 port map( A => ab_2_11_port, B => n3, CI => n31, CO => 
                           CARRYB_2_11_port, S => SUMB_2_11_port);
   S2_2_12 : FA_X1 port map( A => ab_2_12_port, B => n2, CI => n32, CO => 
                           CARRYB_2_12_port, S => SUMB_2_12_port);
   S2_2_13 : FA_X1 port map( A => ab_2_13_port, B => n4, CI => n33, CO => 
                           CARRYB_2_13_port, S => SUMB_2_13_port);
   S2_2_14 : FA_X1 port map( A => ab_2_14_port, B => n5, CI => n47, CO => 
                           CARRYB_2_14_port, S => SUMB_2_14_port);
   S2_2_15 : FA_X1 port map( A => ab_2_15_port, B => n19, CI => n46, CO => 
                           CARRYB_2_15_port, S => SUMB_2_15_port);
   S2_2_16 : FA_X1 port map( A => ab_2_16_port, B => n18, CI => n45, CO => 
                           CARRYB_2_16_port, S => SUMB_2_16_port);
   S2_2_17 : FA_X1 port map( A => ab_2_17_port, B => n17, CI => n44, CO => 
                           CARRYB_2_17_port, S => SUMB_2_17_port);
   S2_2_18 : FA_X1 port map( A => ab_2_18_port, B => n16, CI => n43, CO => 
                           CARRYB_2_18_port, S => SUMB_2_18_port);
   S2_2_19 : FA_X1 port map( A => ab_2_19_port, B => n15, CI => n42, CO => 
                           CARRYB_2_19_port, S => SUMB_2_19_port);
   S2_2_20 : FA_X1 port map( A => ab_2_20_port, B => n14, CI => n41, CO => 
                           CARRYB_2_20_port, S => SUMB_2_20_port);
   S2_2_21 : FA_X1 port map( A => ab_2_21_port, B => n13, CI => n40, CO => 
                           CARRYB_2_21_port, S => SUMB_2_21_port);
   S2_2_22 : FA_X1 port map( A => ab_2_22_port, B => n12, CI => n39, CO => 
                           CARRYB_2_22_port, S => SUMB_2_22_port);
   S2_2_23 : FA_X1 port map( A => ab_2_23_port, B => n11, CI => n38, CO => 
                           CARRYB_2_23_port, S => SUMB_2_23_port);
   S2_2_24 : FA_X1 port map( A => ab_2_24_port, B => n10, CI => n37, CO => 
                           CARRYB_2_24_port, S => SUMB_2_24_port);
   S2_2_25 : FA_X1 port map( A => ab_2_25_port, B => n9, CI => n36, CO => 
                           CARRYB_2_25_port, S => SUMB_2_25_port);
   S2_2_26 : FA_X1 port map( A => ab_2_26_port, B => n8, CI => n35, CO => 
                           CARRYB_2_26_port, S => SUMB_2_26_port);
   S2_2_27 : FA_X1 port map( A => ab_2_27_port, B => n7, CI => n34, CO => 
                           CARRYB_2_27_port, S => SUMB_2_27_port);
   S2_2_28 : FA_X1 port map( A => ab_2_28_port, B => n6, CI => n48, CO => 
                           CARRYB_2_28_port, S => SUMB_2_28_port);
   S2_2_29 : FA_X1 port map( A => ab_2_29_port, B => n61, CI => n62, CO => 
                           n_1062, S => SUMB_2_29_port);
   U2 : AND2_X1 port map( A1 => ab_0_13_port, A2 => ab_1_12_port, ZN => n2);
   U3 : AND2_X1 port map( A1 => ab_0_12_port, A2 => ab_1_11_port, ZN => n3);
   U4 : AND2_X1 port map( A1 => ab_0_14_port, A2 => ab_1_13_port, ZN => n4);
   U5 : AND2_X1 port map( A1 => ab_0_15_port, A2 => ab_1_14_port, ZN => n5);
   U6 : AND2_X1 port map( A1 => ab_0_29_port, A2 => ab_1_28_port, ZN => n6);
   U7 : AND2_X1 port map( A1 => ab_0_28_port, A2 => ab_1_27_port, ZN => n7);
   U8 : AND2_X1 port map( A1 => ab_0_27_port, A2 => ab_1_26_port, ZN => n8);
   U9 : AND2_X1 port map( A1 => ab_0_26_port, A2 => ab_1_25_port, ZN => n9);
   U10 : AND2_X1 port map( A1 => ab_0_25_port, A2 => ab_1_24_port, ZN => n10);
   U11 : AND2_X1 port map( A1 => ab_0_24_port, A2 => ab_1_23_port, ZN => n11);
   U12 : AND2_X1 port map( A1 => ab_0_23_port, A2 => ab_1_22_port, ZN => n12);
   U13 : AND2_X1 port map( A1 => ab_0_22_port, A2 => ab_1_21_port, ZN => n13);
   U14 : AND2_X1 port map( A1 => ab_0_21_port, A2 => ab_1_20_port, ZN => n14);
   U15 : AND2_X1 port map( A1 => ab_0_20_port, A2 => ab_1_19_port, ZN => n15);
   U16 : AND2_X1 port map( A1 => ab_0_19_port, A2 => ab_1_18_port, ZN => n16);
   U17 : AND2_X1 port map( A1 => ab_0_18_port, A2 => ab_1_17_port, ZN => n17);
   U18 : AND2_X1 port map( A1 => ab_0_17_port, A2 => ab_1_16_port, ZN => n18);
   U19 : AND2_X1 port map( A1 => ab_0_16_port, A2 => ab_1_15_port, ZN => n19);
   U20 : XOR2_X1 port map( A => ab_1_11_port, B => ab_0_12_port, Z => n20);
   U21 : AND2_X1 port map( A1 => ab_0_9_port, A2 => ab_1_8_port, ZN => n21);
   U22 : AND2_X1 port map( A1 => ab_0_10_port, A2 => ab_1_9_port, ZN => n22);
   U23 : AND2_X1 port map( A1 => ab_0_2_port, A2 => ab_1_1_port, ZN => n23);
   U24 : AND2_X1 port map( A1 => ab_0_1_port, A2 => ab_1_0_port, ZN => n24);
   U25 : AND2_X1 port map( A1 => ab_0_8_port, A2 => ab_1_7_port, ZN => n25);
   U26 : AND2_X1 port map( A1 => ab_0_7_port, A2 => ab_1_6_port, ZN => n26);
   U27 : AND2_X1 port map( A1 => ab_0_6_port, A2 => ab_1_5_port, ZN => n27);
   U28 : AND2_X1 port map( A1 => ab_0_5_port, A2 => ab_1_4_port, ZN => n28);
   U29 : AND2_X1 port map( A1 => ab_0_4_port, A2 => ab_1_3_port, ZN => n29);
   U30 : AND2_X1 port map( A1 => ab_0_3_port, A2 => ab_1_2_port, ZN => n30);
   U31 : XOR2_X1 port map( A => ab_1_12_port, B => ab_0_13_port, Z => n31);
   U32 : XOR2_X1 port map( A => ab_1_13_port, B => ab_0_14_port, Z => n32);
   U33 : XOR2_X1 port map( A => ab_1_14_port, B => ab_0_15_port, Z => n33);
   U34 : XOR2_X1 port map( A => ab_1_28_port, B => ab_0_29_port, Z => n34);
   U35 : XOR2_X1 port map( A => ab_1_27_port, B => ab_0_28_port, Z => n35);
   U36 : XOR2_X1 port map( A => ab_1_26_port, B => ab_0_27_port, Z => n36);
   U37 : XOR2_X1 port map( A => ab_1_25_port, B => ab_0_26_port, Z => n37);
   U38 : XOR2_X1 port map( A => ab_1_24_port, B => ab_0_25_port, Z => n38);
   U39 : XOR2_X1 port map( A => ab_1_23_port, B => ab_0_24_port, Z => n39);
   U40 : XOR2_X1 port map( A => ab_1_22_port, B => ab_0_23_port, Z => n40);
   U41 : XOR2_X1 port map( A => ab_1_21_port, B => ab_0_22_port, Z => n41);
   U42 : XOR2_X1 port map( A => ab_1_20_port, B => ab_0_21_port, Z => n42);
   U43 : XOR2_X1 port map( A => ab_1_19_port, B => ab_0_20_port, Z => n43);
   U44 : XOR2_X1 port map( A => ab_1_18_port, B => ab_0_19_port, Z => n44);
   U45 : XOR2_X1 port map( A => ab_1_17_port, B => ab_0_18_port, Z => n45);
   U46 : XOR2_X1 port map( A => ab_1_16_port, B => ab_0_17_port, Z => n46);
   U47 : XOR2_X1 port map( A => ab_1_15_port, B => ab_0_16_port, Z => n47);
   U48 : XOR2_X1 port map( A => ab_1_29_port, B => ab_0_30_port, Z => n48);
   U49 : AND2_X1 port map( A1 => ab_0_11_port, A2 => ab_1_10_port, ZN => n49);
   U50 : XOR2_X1 port map( A => ab_1_8_port, B => ab_0_9_port, Z => n50);
   U51 : XOR2_X1 port map( A => ab_1_9_port, B => ab_0_10_port, Z => n51);
   U52 : XOR2_X1 port map( A => ab_1_10_port, B => ab_0_11_port, Z => n52);
   U53 : XOR2_X1 port map( A => ab_1_1_port, B => ab_0_2_port, Z => n53);
   U54 : XOR2_X1 port map( A => ab_1_7_port, B => ab_0_8_port, Z => n54);
   U55 : XOR2_X1 port map( A => ab_1_6_port, B => ab_0_7_port, Z => n55);
   U56 : XOR2_X1 port map( A => ab_1_5_port, B => ab_0_6_port, Z => n56);
   U57 : XOR2_X1 port map( A => ab_1_4_port, B => ab_0_5_port, Z => n57);
   U58 : XOR2_X1 port map( A => ab_1_3_port, B => ab_0_4_port, Z => n58);
   U59 : XOR2_X1 port map( A => ab_1_2_port, B => ab_0_3_port, Z => n59);
   U60 : XOR2_X1 port map( A => ab_1_0_port, B => ab_0_1_port, Z => PRODUCT(1))
                           ;
   U61 : AND2_X1 port map( A1 => ab_0_30_port, A2 => ab_1_29_port, ZN => n61);
   U62 : XOR2_X1 port map( A => ab_0_31_port, B => ab_1_30_port, Z => n62);
   U63 : BUF_X1 port map( A => n144, Z => n86);
   U64 : BUF_X1 port map( A => n143, Z => n82);
   U65 : BUF_X1 port map( A => n144, Z => n85);
   U66 : BUF_X1 port map( A => n143, Z => n83);
   U67 : BUF_X1 port map( A => n142, Z => n80);
   U68 : BUF_X1 port map( A => n141, Z => n77);
   U69 : BUF_X1 port map( A => n142, Z => n79);
   U70 : BUF_X1 port map( A => n144, Z => n87);
   U71 : BUF_X1 port map( A => n168, Z => n89);
   U72 : BUF_X1 port map( A => n169, Z => n91);
   U73 : BUF_X1 port map( A => n170, Z => n93);
   U74 : BUF_X1 port map( A => n171, Z => n96);
   U75 : BUF_X1 port map( A => n172, Z => n99);
   U76 : BUF_X1 port map( A => n173, Z => n102);
   U77 : BUF_X1 port map( A => n174, Z => n105);
   U78 : BUF_X1 port map( A => n175, Z => n108);
   U79 : BUF_X1 port map( A => n176, Z => n111);
   U80 : BUF_X1 port map( A => n168, Z => n88);
   U81 : BUF_X1 port map( A => n169, Z => n90);
   U82 : BUF_X1 port map( A => n170, Z => n92);
   U83 : BUF_X1 port map( A => n172, Z => n98);
   U84 : BUF_X1 port map( A => n171, Z => n95);
   U85 : BUF_X1 port map( A => n174, Z => n104);
   U86 : BUF_X1 port map( A => n175, Z => n107);
   U87 : BUF_X1 port map( A => n173, Z => n101);
   U88 : BUF_X1 port map( A => n176, Z => n110);
   U89 : BUF_X1 port map( A => n136, Z => n64);
   U90 : BUF_X1 port map( A => n136, Z => n63);
   U91 : BUF_X1 port map( A => n137, Z => n66);
   U92 : BUF_X1 port map( A => n137, Z => n65);
   U93 : BUF_X1 port map( A => n141, Z => n76);
   U94 : BUF_X1 port map( A => n140, Z => n74);
   U95 : BUF_X1 port map( A => n140, Z => n73);
   U96 : BUF_X1 port map( A => n139, Z => n71);
   U97 : BUF_X1 port map( A => n139, Z => n70);
   U98 : BUF_X1 port map( A => n138, Z => n68);
   U99 : BUF_X1 port map( A => n138, Z => n67);
   U100 : BUF_X1 port map( A => n175, Z => n109);
   U101 : BUF_X1 port map( A => n143, Z => n84);
   U102 : BUF_X1 port map( A => n174, Z => n106);
   U103 : BUF_X1 port map( A => n142, Z => n81);
   U104 : BUF_X1 port map( A => n173, Z => n103);
   U105 : BUF_X1 port map( A => n141, Z => n78);
   U106 : BUF_X1 port map( A => n172, Z => n100);
   U107 : BUF_X1 port map( A => n140, Z => n75);
   U108 : BUF_X1 port map( A => n171, Z => n97);
   U109 : BUF_X1 port map( A => n139, Z => n72);
   U110 : BUF_X1 port map( A => n170, Z => n94);
   U111 : BUF_X1 port map( A => n138, Z => n69);
   U112 : BUF_X1 port map( A => n176, Z => n112);
   U113 : INV_X1 port map( A => B(13), ZN => n163);
   U114 : INV_X1 port map( A => B(14), ZN => n162);
   U115 : INV_X1 port map( A => B(15), ZN => n161);
   U116 : INV_X1 port map( A => B(16), ZN => n160);
   U117 : INV_X1 port map( A => B(17), ZN => n159);
   U118 : INV_X1 port map( A => B(18), ZN => n158);
   U119 : INV_X1 port map( A => B(19), ZN => n157);
   U120 : INV_X1 port map( A => B(20), ZN => n156);
   U121 : INV_X1 port map( A => B(21), ZN => n155);
   U122 : INV_X1 port map( A => B(12), ZN => n164);
   U123 : INV_X1 port map( A => B(22), ZN => n154);
   U124 : INV_X1 port map( A => B(23), ZN => n153);
   U125 : INV_X1 port map( A => B(24), ZN => n152);
   U126 : INV_X1 port map( A => B(25), ZN => n151);
   U127 : INV_X1 port map( A => B(26), ZN => n150);
   U128 : INV_X1 port map( A => A(31), ZN => n113);
   U129 : INV_X1 port map( A => B(27), ZN => n149);
   U130 : INV_X1 port map( A => B(28), ZN => n148);
   U131 : INV_X1 port map( A => B(29), ZN => n147);
   U132 : INV_X1 port map( A => A(1), ZN => n143);
   U133 : INV_X1 port map( A => A(0), ZN => n144);
   U134 : INV_X1 port map( A => A(2), ZN => n142);
   U135 : INV_X1 port map( A => A(3), ZN => n141);
   U136 : INV_X1 port map( A => B(30), ZN => n146);
   U137 : INV_X1 port map( A => B(31), ZN => n145);
   U138 : INV_X1 port map( A => A(9), ZN => n135);
   U139 : INV_X1 port map( A => B(9), ZN => n167);
   U140 : INV_X1 port map( A => B(10), ZN => n166);
   U141 : INV_X1 port map( A => A(10), ZN => n134);
   U142 : INV_X1 port map( A => B(11), ZN => n165);
   U143 : INV_X1 port map( A => A(11), ZN => n133);
   U144 : INV_X1 port map( A => B(6), ZN => n170);
   U145 : INV_X1 port map( A => B(5), ZN => n171);
   U146 : INV_X1 port map( A => B(4), ZN => n172);
   U147 : INV_X1 port map( A => B(3), ZN => n173);
   U148 : INV_X1 port map( A => B(2), ZN => n174);
   U149 : INV_X1 port map( A => A(4), ZN => n140);
   U150 : INV_X1 port map( A => A(5), ZN => n139);
   U151 : INV_X1 port map( A => A(6), ZN => n138);
   U152 : INV_X1 port map( A => B(1), ZN => n175);
   U153 : INV_X1 port map( A => B(0), ZN => n176);
   U154 : INV_X1 port map( A => A(7), ZN => n137);
   U155 : INV_X1 port map( A => B(7), ZN => n169);
   U156 : INV_X1 port map( A => B(8), ZN => n168);
   U157 : INV_X1 port map( A => A(8), ZN => n136);
   U158 : INV_X1 port map( A => A(13), ZN => n131);
   U159 : INV_X1 port map( A => A(14), ZN => n130);
   U160 : INV_X1 port map( A => A(15), ZN => n129);
   U161 : INV_X1 port map( A => A(16), ZN => n128);
   U162 : INV_X1 port map( A => A(17), ZN => n127);
   U163 : INV_X1 port map( A => A(18), ZN => n126);
   U164 : INV_X1 port map( A => A(12), ZN => n132);
   U165 : INV_X1 port map( A => A(19), ZN => n125);
   U166 : INV_X1 port map( A => A(20), ZN => n124);
   U167 : INV_X1 port map( A => A(21), ZN => n123);
   U168 : INV_X1 port map( A => A(22), ZN => n122);
   U169 : INV_X1 port map( A => A(23), ZN => n121);
   U170 : INV_X1 port map( A => A(24), ZN => n120);
   U171 : INV_X1 port map( A => A(25), ZN => n119);
   U172 : INV_X1 port map( A => A(26), ZN => n118);
   U173 : INV_X1 port map( A => A(27), ZN => n117);
   U174 : INV_X1 port map( A => A(28), ZN => n116);
   U175 : INV_X1 port map( A => A(29), ZN => n115);
   U176 : INV_X1 port map( A => A(30), ZN => n114);
   U177 : NOR2_X1 port map( A1 => n135, A2 => n167, ZN => ab_9_9_port);
   U178 : NOR2_X1 port map( A1 => n135, A2 => n88, ZN => ab_9_8_port);
   U179 : NOR2_X1 port map( A1 => n135, A2 => n90, ZN => ab_9_7_port);
   U180 : NOR2_X1 port map( A1 => n135, A2 => n92, ZN => ab_9_6_port);
   U181 : NOR2_X1 port map( A1 => n135, A2 => n95, ZN => ab_9_5_port);
   U182 : NOR2_X1 port map( A1 => n135, A2 => n98, ZN => ab_9_4_port);
   U183 : NOR2_X1 port map( A1 => n135, A2 => n101, ZN => ab_9_3_port);
   U184 : NOR2_X1 port map( A1 => n135, A2 => n104, ZN => ab_9_2_port);
   U185 : NOR2_X1 port map( A1 => n135, A2 => n154, ZN => ab_9_22_port);
   U186 : NOR2_X1 port map( A1 => n135, A2 => n155, ZN => ab_9_21_port);
   U187 : NOR2_X1 port map( A1 => n135, A2 => n156, ZN => ab_9_20_port);
   U188 : NOR2_X1 port map( A1 => n135, A2 => n107, ZN => ab_9_1_port);
   U189 : NOR2_X1 port map( A1 => n135, A2 => n157, ZN => ab_9_19_port);
   U190 : NOR2_X1 port map( A1 => n135, A2 => n158, ZN => ab_9_18_port);
   U191 : NOR2_X1 port map( A1 => n135, A2 => n159, ZN => ab_9_17_port);
   U192 : NOR2_X1 port map( A1 => n135, A2 => n160, ZN => ab_9_16_port);
   U193 : NOR2_X1 port map( A1 => n135, A2 => n161, ZN => ab_9_15_port);
   U194 : NOR2_X1 port map( A1 => n135, A2 => n162, ZN => ab_9_14_port);
   U195 : NOR2_X1 port map( A1 => n135, A2 => n163, ZN => ab_9_13_port);
   U196 : NOR2_X1 port map( A1 => n135, A2 => n164, ZN => ab_9_12_port);
   U197 : NOR2_X1 port map( A1 => n135, A2 => n165, ZN => ab_9_11_port);
   U198 : NOR2_X1 port map( A1 => n135, A2 => n166, ZN => ab_9_10_port);
   U199 : NOR2_X1 port map( A1 => n135, A2 => n110, ZN => ab_9_0_port);
   U200 : NOR2_X1 port map( A1 => n167, A2 => n64, ZN => ab_8_9_port);
   U201 : NOR2_X1 port map( A1 => n88, A2 => n64, ZN => ab_8_8_port);
   U202 : NOR2_X1 port map( A1 => n90, A2 => n64, ZN => ab_8_7_port);
   U203 : NOR2_X1 port map( A1 => n92, A2 => n64, ZN => ab_8_6_port);
   U204 : NOR2_X1 port map( A1 => n95, A2 => n64, ZN => ab_8_5_port);
   U205 : NOR2_X1 port map( A1 => n98, A2 => n64, ZN => ab_8_4_port);
   U206 : NOR2_X1 port map( A1 => n101, A2 => n64, ZN => ab_8_3_port);
   U207 : NOR2_X1 port map( A1 => n104, A2 => n64, ZN => ab_8_2_port);
   U208 : NOR2_X1 port map( A1 => n153, A2 => n64, ZN => ab_8_23_port);
   U209 : NOR2_X1 port map( A1 => n154, A2 => n64, ZN => ab_8_22_port);
   U210 : NOR2_X1 port map( A1 => n155, A2 => n64, ZN => ab_8_21_port);
   U211 : NOR2_X1 port map( A1 => n156, A2 => n64, ZN => ab_8_20_port);
   U212 : NOR2_X1 port map( A1 => n107, A2 => n63, ZN => ab_8_1_port);
   U213 : NOR2_X1 port map( A1 => n157, A2 => n63, ZN => ab_8_19_port);
   U214 : NOR2_X1 port map( A1 => n158, A2 => n63, ZN => ab_8_18_port);
   U215 : NOR2_X1 port map( A1 => n159, A2 => n63, ZN => ab_8_17_port);
   U216 : NOR2_X1 port map( A1 => n160, A2 => n63, ZN => ab_8_16_port);
   U217 : NOR2_X1 port map( A1 => n161, A2 => n63, ZN => ab_8_15_port);
   U218 : NOR2_X1 port map( A1 => n162, A2 => n63, ZN => ab_8_14_port);
   U219 : NOR2_X1 port map( A1 => n163, A2 => n63, ZN => ab_8_13_port);
   U220 : NOR2_X1 port map( A1 => n164, A2 => n63, ZN => ab_8_12_port);
   U221 : NOR2_X1 port map( A1 => n165, A2 => n63, ZN => ab_8_11_port);
   U222 : NOR2_X1 port map( A1 => n166, A2 => n63, ZN => ab_8_10_port);
   U223 : NOR2_X1 port map( A1 => n110, A2 => n63, ZN => ab_8_0_port);
   U224 : NOR2_X1 port map( A1 => n167, A2 => n65, ZN => ab_7_9_port);
   U225 : NOR2_X1 port map( A1 => n88, A2 => n66, ZN => ab_7_8_port);
   U226 : NOR2_X1 port map( A1 => n90, A2 => n66, ZN => ab_7_7_port);
   U227 : NOR2_X1 port map( A1 => n92, A2 => n66, ZN => ab_7_6_port);
   U228 : NOR2_X1 port map( A1 => n95, A2 => n66, ZN => ab_7_5_port);
   U229 : NOR2_X1 port map( A1 => n98, A2 => n66, ZN => ab_7_4_port);
   U230 : NOR2_X1 port map( A1 => n101, A2 => n66, ZN => ab_7_3_port);
   U231 : NOR2_X1 port map( A1 => n104, A2 => n66, ZN => ab_7_2_port);
   U232 : NOR2_X1 port map( A1 => n152, A2 => n66, ZN => ab_7_24_port);
   U233 : NOR2_X1 port map( A1 => n153, A2 => n66, ZN => ab_7_23_port);
   U234 : NOR2_X1 port map( A1 => n154, A2 => n66, ZN => ab_7_22_port);
   U235 : NOR2_X1 port map( A1 => n155, A2 => n66, ZN => ab_7_21_port);
   U236 : NOR2_X1 port map( A1 => n156, A2 => n66, ZN => ab_7_20_port);
   U237 : NOR2_X1 port map( A1 => n107, A2 => n65, ZN => ab_7_1_port);
   U238 : NOR2_X1 port map( A1 => n157, A2 => n65, ZN => ab_7_19_port);
   U239 : NOR2_X1 port map( A1 => n158, A2 => n65, ZN => ab_7_18_port);
   U240 : NOR2_X1 port map( A1 => n159, A2 => n65, ZN => ab_7_17_port);
   U241 : NOR2_X1 port map( A1 => n160, A2 => n65, ZN => ab_7_16_port);
   U242 : NOR2_X1 port map( A1 => n161, A2 => n65, ZN => ab_7_15_port);
   U243 : NOR2_X1 port map( A1 => n162, A2 => n65, ZN => ab_7_14_port);
   U244 : NOR2_X1 port map( A1 => n163, A2 => n65, ZN => ab_7_13_port);
   U245 : NOR2_X1 port map( A1 => n164, A2 => n65, ZN => ab_7_12_port);
   U246 : NOR2_X1 port map( A1 => n165, A2 => n65, ZN => ab_7_11_port);
   U247 : NOR2_X1 port map( A1 => n166, A2 => n65, ZN => ab_7_10_port);
   U248 : NOR2_X1 port map( A1 => n110, A2 => n65, ZN => ab_7_0_port);
   U249 : NOR2_X1 port map( A1 => n167, A2 => n69, ZN => ab_6_9_port);
   U250 : NOR2_X1 port map( A1 => n88, A2 => n69, ZN => ab_6_8_port);
   U251 : NOR2_X1 port map( A1 => n90, A2 => n68, ZN => ab_6_7_port);
   U252 : NOR2_X1 port map( A1 => n92, A2 => n68, ZN => ab_6_6_port);
   U253 : NOR2_X1 port map( A1 => n95, A2 => n68, ZN => ab_6_5_port);
   U254 : NOR2_X1 port map( A1 => n98, A2 => n68, ZN => ab_6_4_port);
   U255 : NOR2_X1 port map( A1 => n101, A2 => n68, ZN => ab_6_3_port);
   U256 : NOR2_X1 port map( A1 => n104, A2 => n68, ZN => ab_6_2_port);
   U257 : NOR2_X1 port map( A1 => n151, A2 => n68, ZN => ab_6_25_port);
   U258 : NOR2_X1 port map( A1 => n152, A2 => n68, ZN => ab_6_24_port);
   U259 : NOR2_X1 port map( A1 => n153, A2 => n68, ZN => ab_6_23_port);
   U260 : NOR2_X1 port map( A1 => n154, A2 => n68, ZN => ab_6_22_port);
   U261 : NOR2_X1 port map( A1 => n155, A2 => n68, ZN => ab_6_21_port);
   U262 : NOR2_X1 port map( A1 => n156, A2 => n68, ZN => ab_6_20_port);
   U263 : NOR2_X1 port map( A1 => n107, A2 => n67, ZN => ab_6_1_port);
   U264 : NOR2_X1 port map( A1 => n157, A2 => n67, ZN => ab_6_19_port);
   U265 : NOR2_X1 port map( A1 => n158, A2 => n67, ZN => ab_6_18_port);
   U266 : NOR2_X1 port map( A1 => n159, A2 => n67, ZN => ab_6_17_port);
   U267 : NOR2_X1 port map( A1 => n160, A2 => n67, ZN => ab_6_16_port);
   U268 : NOR2_X1 port map( A1 => n161, A2 => n67, ZN => ab_6_15_port);
   U269 : NOR2_X1 port map( A1 => n162, A2 => n67, ZN => ab_6_14_port);
   U270 : NOR2_X1 port map( A1 => n163, A2 => n67, ZN => ab_6_13_port);
   U271 : NOR2_X1 port map( A1 => n164, A2 => n67, ZN => ab_6_12_port);
   U272 : NOR2_X1 port map( A1 => n165, A2 => n67, ZN => ab_6_11_port);
   U273 : NOR2_X1 port map( A1 => n166, A2 => n67, ZN => ab_6_10_port);
   U274 : NOR2_X1 port map( A1 => n110, A2 => n67, ZN => ab_6_0_port);
   U275 : NOR2_X1 port map( A1 => n167, A2 => n72, ZN => ab_5_9_port);
   U276 : NOR2_X1 port map( A1 => n88, A2 => n72, ZN => ab_5_8_port);
   U277 : NOR2_X1 port map( A1 => n90, A2 => n72, ZN => ab_5_7_port);
   U278 : NOR2_X1 port map( A1 => n92, A2 => n71, ZN => ab_5_6_port);
   U279 : NOR2_X1 port map( A1 => n95, A2 => n71, ZN => ab_5_5_port);
   U280 : NOR2_X1 port map( A1 => n98, A2 => n71, ZN => ab_5_4_port);
   U281 : NOR2_X1 port map( A1 => n101, A2 => n71, ZN => ab_5_3_port);
   U282 : NOR2_X1 port map( A1 => n104, A2 => n71, ZN => ab_5_2_port);
   U283 : NOR2_X1 port map( A1 => n150, A2 => n71, ZN => ab_5_26_port);
   U284 : NOR2_X1 port map( A1 => n151, A2 => n71, ZN => ab_5_25_port);
   U285 : NOR2_X1 port map( A1 => n152, A2 => n71, ZN => ab_5_24_port);
   U286 : NOR2_X1 port map( A1 => n153, A2 => n71, ZN => ab_5_23_port);
   U287 : NOR2_X1 port map( A1 => n154, A2 => n71, ZN => ab_5_22_port);
   U288 : NOR2_X1 port map( A1 => n155, A2 => n71, ZN => ab_5_21_port);
   U289 : NOR2_X1 port map( A1 => n156, A2 => n71, ZN => ab_5_20_port);
   U290 : NOR2_X1 port map( A1 => n107, A2 => n70, ZN => ab_5_1_port);
   U291 : NOR2_X1 port map( A1 => n157, A2 => n70, ZN => ab_5_19_port);
   U292 : NOR2_X1 port map( A1 => n158, A2 => n70, ZN => ab_5_18_port);
   U293 : NOR2_X1 port map( A1 => n159, A2 => n70, ZN => ab_5_17_port);
   U294 : NOR2_X1 port map( A1 => n160, A2 => n70, ZN => ab_5_16_port);
   U295 : NOR2_X1 port map( A1 => n161, A2 => n70, ZN => ab_5_15_port);
   U296 : NOR2_X1 port map( A1 => n162, A2 => n70, ZN => ab_5_14_port);
   U297 : NOR2_X1 port map( A1 => n163, A2 => n70, ZN => ab_5_13_port);
   U298 : NOR2_X1 port map( A1 => n164, A2 => n70, ZN => ab_5_12_port);
   U299 : NOR2_X1 port map( A1 => n165, A2 => n70, ZN => ab_5_11_port);
   U300 : NOR2_X1 port map( A1 => n166, A2 => n70, ZN => ab_5_10_port);
   U301 : NOR2_X1 port map( A1 => n110, A2 => n70, ZN => ab_5_0_port);
   U302 : NOR2_X1 port map( A1 => n167, A2 => n75, ZN => ab_4_9_port);
   U303 : NOR2_X1 port map( A1 => n88, A2 => n75, ZN => ab_4_8_port);
   U304 : NOR2_X1 port map( A1 => n90, A2 => n75, ZN => ab_4_7_port);
   U305 : NOR2_X1 port map( A1 => n92, A2 => n75, ZN => ab_4_6_port);
   U306 : NOR2_X1 port map( A1 => n95, A2 => n74, ZN => ab_4_5_port);
   U307 : NOR2_X1 port map( A1 => n98, A2 => n74, ZN => ab_4_4_port);
   U308 : NOR2_X1 port map( A1 => n101, A2 => n74, ZN => ab_4_3_port);
   U309 : NOR2_X1 port map( A1 => n104, A2 => n74, ZN => ab_4_2_port);
   U310 : NOR2_X1 port map( A1 => n149, A2 => n74, ZN => ab_4_27_port);
   U311 : NOR2_X1 port map( A1 => n150, A2 => n74, ZN => ab_4_26_port);
   U312 : NOR2_X1 port map( A1 => n151, A2 => n74, ZN => ab_4_25_port);
   U313 : NOR2_X1 port map( A1 => n152, A2 => n74, ZN => ab_4_24_port);
   U314 : NOR2_X1 port map( A1 => n153, A2 => n74, ZN => ab_4_23_port);
   U315 : NOR2_X1 port map( A1 => n154, A2 => n74, ZN => ab_4_22_port);
   U316 : NOR2_X1 port map( A1 => n155, A2 => n74, ZN => ab_4_21_port);
   U317 : NOR2_X1 port map( A1 => n156, A2 => n74, ZN => ab_4_20_port);
   U318 : NOR2_X1 port map( A1 => n107, A2 => n73, ZN => ab_4_1_port);
   U319 : NOR2_X1 port map( A1 => n157, A2 => n73, ZN => ab_4_19_port);
   U320 : NOR2_X1 port map( A1 => n158, A2 => n73, ZN => ab_4_18_port);
   U321 : NOR2_X1 port map( A1 => n159, A2 => n73, ZN => ab_4_17_port);
   U322 : NOR2_X1 port map( A1 => n160, A2 => n73, ZN => ab_4_16_port);
   U323 : NOR2_X1 port map( A1 => n161, A2 => n73, ZN => ab_4_15_port);
   U324 : NOR2_X1 port map( A1 => n162, A2 => n73, ZN => ab_4_14_port);
   U325 : NOR2_X1 port map( A1 => n163, A2 => n73, ZN => ab_4_13_port);
   U326 : NOR2_X1 port map( A1 => n164, A2 => n73, ZN => ab_4_12_port);
   U327 : NOR2_X1 port map( A1 => n165, A2 => n73, ZN => ab_4_11_port);
   U328 : NOR2_X1 port map( A1 => n166, A2 => n73, ZN => ab_4_10_port);
   U329 : NOR2_X1 port map( A1 => n110, A2 => n73, ZN => ab_4_0_port);
   U330 : NOR2_X1 port map( A1 => n167, A2 => n78, ZN => ab_3_9_port);
   U331 : NOR2_X1 port map( A1 => n88, A2 => n78, ZN => ab_3_8_port);
   U332 : NOR2_X1 port map( A1 => n90, A2 => n78, ZN => ab_3_7_port);
   U333 : NOR2_X1 port map( A1 => n92, A2 => n78, ZN => ab_3_6_port);
   U334 : NOR2_X1 port map( A1 => n95, A2 => n78, ZN => ab_3_5_port);
   U335 : NOR2_X1 port map( A1 => n98, A2 => n77, ZN => ab_3_4_port);
   U336 : NOR2_X1 port map( A1 => n101, A2 => n77, ZN => ab_3_3_port);
   U337 : NOR2_X1 port map( A1 => n104, A2 => n77, ZN => ab_3_2_port);
   U338 : NOR2_X1 port map( A1 => n148, A2 => n77, ZN => ab_3_28_port);
   U339 : NOR2_X1 port map( A1 => n149, A2 => n77, ZN => ab_3_27_port);
   U340 : NOR2_X1 port map( A1 => n150, A2 => n77, ZN => ab_3_26_port);
   U341 : NOR2_X1 port map( A1 => n151, A2 => n77, ZN => ab_3_25_port);
   U342 : NOR2_X1 port map( A1 => n152, A2 => n77, ZN => ab_3_24_port);
   U343 : NOR2_X1 port map( A1 => n153, A2 => n77, ZN => ab_3_23_port);
   U344 : NOR2_X1 port map( A1 => n154, A2 => n77, ZN => ab_3_22_port);
   U345 : NOR2_X1 port map( A1 => n155, A2 => n77, ZN => ab_3_21_port);
   U346 : NOR2_X1 port map( A1 => n156, A2 => n77, ZN => ab_3_20_port);
   U347 : NOR2_X1 port map( A1 => n107, A2 => n76, ZN => ab_3_1_port);
   U348 : NOR2_X1 port map( A1 => n157, A2 => n76, ZN => ab_3_19_port);
   U349 : NOR2_X1 port map( A1 => n158, A2 => n76, ZN => ab_3_18_port);
   U350 : NOR2_X1 port map( A1 => n159, A2 => n76, ZN => ab_3_17_port);
   U351 : NOR2_X1 port map( A1 => n160, A2 => n76, ZN => ab_3_16_port);
   U352 : NOR2_X1 port map( A1 => n161, A2 => n76, ZN => ab_3_15_port);
   U353 : NOR2_X1 port map( A1 => n162, A2 => n76, ZN => ab_3_14_port);
   U354 : NOR2_X1 port map( A1 => n163, A2 => n76, ZN => ab_3_13_port);
   U355 : NOR2_X1 port map( A1 => n164, A2 => n76, ZN => ab_3_12_port);
   U356 : NOR2_X1 port map( A1 => n165, A2 => n76, ZN => ab_3_11_port);
   U357 : NOR2_X1 port map( A1 => n166, A2 => n76, ZN => ab_3_10_port);
   U358 : NOR2_X1 port map( A1 => n110, A2 => n76, ZN => ab_3_0_port);
   U359 : NOR2_X1 port map( A1 => n110, A2 => n113, ZN => ab_31_0_port);
   U360 : NOR2_X1 port map( A1 => n107, A2 => n114, ZN => ab_30_1_port);
   U361 : NOR2_X1 port map( A1 => n110, A2 => n114, ZN => ab_30_0_port);
   U362 : NOR2_X1 port map( A1 => n167, A2 => n81, ZN => ab_2_9_port);
   U363 : NOR2_X1 port map( A1 => n88, A2 => n81, ZN => ab_2_8_port);
   U364 : NOR2_X1 port map( A1 => n90, A2 => n81, ZN => ab_2_7_port);
   U365 : NOR2_X1 port map( A1 => n92, A2 => n81, ZN => ab_2_6_port);
   U366 : NOR2_X1 port map( A1 => n95, A2 => n81, ZN => ab_2_5_port);
   U367 : NOR2_X1 port map( A1 => n98, A2 => n81, ZN => ab_2_4_port);
   U368 : NOR2_X1 port map( A1 => n101, A2 => n80, ZN => ab_2_3_port);
   U369 : NOR2_X1 port map( A1 => n104, A2 => n80, ZN => ab_2_2_port);
   U370 : NOR2_X1 port map( A1 => n147, A2 => n80, ZN => ab_2_29_port);
   U371 : NOR2_X1 port map( A1 => n148, A2 => n80, ZN => ab_2_28_port);
   U372 : NOR2_X1 port map( A1 => n149, A2 => n80, ZN => ab_2_27_port);
   U373 : NOR2_X1 port map( A1 => n150, A2 => n80, ZN => ab_2_26_port);
   U374 : NOR2_X1 port map( A1 => n151, A2 => n80, ZN => ab_2_25_port);
   U375 : NOR2_X1 port map( A1 => n152, A2 => n80, ZN => ab_2_24_port);
   U376 : NOR2_X1 port map( A1 => n153, A2 => n80, ZN => ab_2_23_port);
   U377 : NOR2_X1 port map( A1 => n154, A2 => n80, ZN => ab_2_22_port);
   U378 : NOR2_X1 port map( A1 => n155, A2 => n80, ZN => ab_2_21_port);
   U379 : NOR2_X1 port map( A1 => n156, A2 => n80, ZN => ab_2_20_port);
   U380 : NOR2_X1 port map( A1 => n107, A2 => n79, ZN => ab_2_1_port);
   U381 : NOR2_X1 port map( A1 => n157, A2 => n79, ZN => ab_2_19_port);
   U382 : NOR2_X1 port map( A1 => n158, A2 => n79, ZN => ab_2_18_port);
   U383 : NOR2_X1 port map( A1 => n159, A2 => n79, ZN => ab_2_17_port);
   U384 : NOR2_X1 port map( A1 => n160, A2 => n79, ZN => ab_2_16_port);
   U385 : NOR2_X1 port map( A1 => n161, A2 => n79, ZN => ab_2_15_port);
   U386 : NOR2_X1 port map( A1 => n162, A2 => n79, ZN => ab_2_14_port);
   U387 : NOR2_X1 port map( A1 => n163, A2 => n79, ZN => ab_2_13_port);
   U388 : NOR2_X1 port map( A1 => n164, A2 => n79, ZN => ab_2_12_port);
   U389 : NOR2_X1 port map( A1 => n165, A2 => n79, ZN => ab_2_11_port);
   U390 : NOR2_X1 port map( A1 => n166, A2 => n79, ZN => ab_2_10_port);
   U391 : NOR2_X1 port map( A1 => n110, A2 => n79, ZN => ab_2_0_port);
   U392 : NOR2_X1 port map( A1 => n104, A2 => n115, ZN => ab_29_2_port);
   U393 : NOR2_X1 port map( A1 => n107, A2 => n115, ZN => ab_29_1_port);
   U394 : NOR2_X1 port map( A1 => n110, A2 => n115, ZN => ab_29_0_port);
   U395 : NOR2_X1 port map( A1 => n101, A2 => n116, ZN => ab_28_3_port);
   U396 : NOR2_X1 port map( A1 => n104, A2 => n116, ZN => ab_28_2_port);
   U397 : NOR2_X1 port map( A1 => n107, A2 => n116, ZN => ab_28_1_port);
   U398 : NOR2_X1 port map( A1 => n110, A2 => n116, ZN => ab_28_0_port);
   U399 : NOR2_X1 port map( A1 => n98, A2 => n117, ZN => ab_27_4_port);
   U400 : NOR2_X1 port map( A1 => n101, A2 => n117, ZN => ab_27_3_port);
   U401 : NOR2_X1 port map( A1 => n104, A2 => n117, ZN => ab_27_2_port);
   U402 : NOR2_X1 port map( A1 => n107, A2 => n117, ZN => ab_27_1_port);
   U403 : NOR2_X1 port map( A1 => n111, A2 => n117, ZN => ab_27_0_port);
   U404 : NOR2_X1 port map( A1 => n95, A2 => n118, ZN => ab_26_5_port);
   U405 : NOR2_X1 port map( A1 => n98, A2 => n118, ZN => ab_26_4_port);
   U406 : NOR2_X1 port map( A1 => n101, A2 => n118, ZN => ab_26_3_port);
   U407 : NOR2_X1 port map( A1 => n104, A2 => n118, ZN => ab_26_2_port);
   U408 : NOR2_X1 port map( A1 => n108, A2 => n118, ZN => ab_26_1_port);
   U409 : NOR2_X1 port map( A1 => n111, A2 => n118, ZN => ab_26_0_port);
   U410 : NOR2_X1 port map( A1 => n92, A2 => n119, ZN => ab_25_6_port);
   U411 : NOR2_X1 port map( A1 => n95, A2 => n119, ZN => ab_25_5_port);
   U412 : NOR2_X1 port map( A1 => n98, A2 => n119, ZN => ab_25_4_port);
   U413 : NOR2_X1 port map( A1 => n101, A2 => n119, ZN => ab_25_3_port);
   U414 : NOR2_X1 port map( A1 => n105, A2 => n119, ZN => ab_25_2_port);
   U415 : NOR2_X1 port map( A1 => n108, A2 => n119, ZN => ab_25_1_port);
   U416 : NOR2_X1 port map( A1 => n111, A2 => n119, ZN => ab_25_0_port);
   U417 : NOR2_X1 port map( A1 => n90, A2 => n120, ZN => ab_24_7_port);
   U418 : NOR2_X1 port map( A1 => n92, A2 => n120, ZN => ab_24_6_port);
   U419 : NOR2_X1 port map( A1 => n95, A2 => n120, ZN => ab_24_5_port);
   U420 : NOR2_X1 port map( A1 => n98, A2 => n120, ZN => ab_24_4_port);
   U421 : NOR2_X1 port map( A1 => n102, A2 => n120, ZN => ab_24_3_port);
   U422 : NOR2_X1 port map( A1 => n105, A2 => n120, ZN => ab_24_2_port);
   U423 : NOR2_X1 port map( A1 => n108, A2 => n120, ZN => ab_24_1_port);
   U424 : NOR2_X1 port map( A1 => n111, A2 => n120, ZN => ab_24_0_port);
   U425 : NOR2_X1 port map( A1 => n88, A2 => n121, ZN => ab_23_8_port);
   U426 : NOR2_X1 port map( A1 => n90, A2 => n121, ZN => ab_23_7_port);
   U427 : NOR2_X1 port map( A1 => n92, A2 => n121, ZN => ab_23_6_port);
   U428 : NOR2_X1 port map( A1 => n95, A2 => n121, ZN => ab_23_5_port);
   U429 : NOR2_X1 port map( A1 => n99, A2 => n121, ZN => ab_23_4_port);
   U430 : NOR2_X1 port map( A1 => n102, A2 => n121, ZN => ab_23_3_port);
   U431 : NOR2_X1 port map( A1 => n105, A2 => n121, ZN => ab_23_2_port);
   U432 : NOR2_X1 port map( A1 => n108, A2 => n121, ZN => ab_23_1_port);
   U433 : NOR2_X1 port map( A1 => n111, A2 => n121, ZN => ab_23_0_port);
   U434 : NOR2_X1 port map( A1 => n167, A2 => n122, ZN => ab_22_9_port);
   U435 : NOR2_X1 port map( A1 => n88, A2 => n122, ZN => ab_22_8_port);
   U436 : NOR2_X1 port map( A1 => n90, A2 => n122, ZN => ab_22_7_port);
   U437 : NOR2_X1 port map( A1 => n92, A2 => n122, ZN => ab_22_6_port);
   U438 : NOR2_X1 port map( A1 => n96, A2 => n122, ZN => ab_22_5_port);
   U439 : NOR2_X1 port map( A1 => n99, A2 => n122, ZN => ab_22_4_port);
   U440 : NOR2_X1 port map( A1 => n102, A2 => n122, ZN => ab_22_3_port);
   U441 : NOR2_X1 port map( A1 => n105, A2 => n122, ZN => ab_22_2_port);
   U442 : NOR2_X1 port map( A1 => n108, A2 => n122, ZN => ab_22_1_port);
   U443 : NOR2_X1 port map( A1 => n111, A2 => n122, ZN => ab_22_0_port);
   U444 : NOR2_X1 port map( A1 => n167, A2 => n123, ZN => ab_21_9_port);
   U445 : NOR2_X1 port map( A1 => n88, A2 => n123, ZN => ab_21_8_port);
   U446 : NOR2_X1 port map( A1 => n90, A2 => n123, ZN => ab_21_7_port);
   U447 : NOR2_X1 port map( A1 => n93, A2 => n123, ZN => ab_21_6_port);
   U448 : NOR2_X1 port map( A1 => n96, A2 => n123, ZN => ab_21_5_port);
   U449 : NOR2_X1 port map( A1 => n99, A2 => n123, ZN => ab_21_4_port);
   U450 : NOR2_X1 port map( A1 => n102, A2 => n123, ZN => ab_21_3_port);
   U451 : NOR2_X1 port map( A1 => n105, A2 => n123, ZN => ab_21_2_port);
   U452 : NOR2_X1 port map( A1 => n108, A2 => n123, ZN => ab_21_1_port);
   U453 : NOR2_X1 port map( A1 => n166, A2 => n123, ZN => ab_21_10_port);
   U454 : NOR2_X1 port map( A1 => n111, A2 => n123, ZN => ab_21_0_port);
   U455 : NOR2_X1 port map( A1 => n167, A2 => n124, ZN => ab_20_9_port);
   U456 : NOR2_X1 port map( A1 => n88, A2 => n124, ZN => ab_20_8_port);
   U457 : NOR2_X1 port map( A1 => n91, A2 => n124, ZN => ab_20_7_port);
   U458 : NOR2_X1 port map( A1 => n93, A2 => n124, ZN => ab_20_6_port);
   U459 : NOR2_X1 port map( A1 => n96, A2 => n124, ZN => ab_20_5_port);
   U460 : NOR2_X1 port map( A1 => n99, A2 => n124, ZN => ab_20_4_port);
   U461 : NOR2_X1 port map( A1 => n102, A2 => n124, ZN => ab_20_3_port);
   U462 : NOR2_X1 port map( A1 => n105, A2 => n124, ZN => ab_20_2_port);
   U463 : NOR2_X1 port map( A1 => n108, A2 => n124, ZN => ab_20_1_port);
   U464 : NOR2_X1 port map( A1 => n165, A2 => n124, ZN => ab_20_11_port);
   U465 : NOR2_X1 port map( A1 => n166, A2 => n124, ZN => ab_20_10_port);
   U466 : NOR2_X1 port map( A1 => n111, A2 => n124, ZN => ab_20_0_port);
   U467 : NOR2_X1 port map( A1 => n167, A2 => n84, ZN => ab_1_9_port);
   U468 : NOR2_X1 port map( A1 => n89, A2 => n84, ZN => ab_1_8_port);
   U469 : NOR2_X1 port map( A1 => n91, A2 => n84, ZN => ab_1_7_port);
   U470 : NOR2_X1 port map( A1 => n93, A2 => n84, ZN => ab_1_6_port);
   U471 : NOR2_X1 port map( A1 => n96, A2 => n84, ZN => ab_1_5_port);
   U472 : NOR2_X1 port map( A1 => n99, A2 => n84, ZN => ab_1_4_port);
   U473 : NOR2_X1 port map( A1 => n102, A2 => n84, ZN => ab_1_3_port);
   U474 : NOR2_X1 port map( A1 => n146, A2 => n83, ZN => ab_1_30_port);
   U475 : NOR2_X1 port map( A1 => n105, A2 => n83, ZN => ab_1_2_port);
   U476 : NOR2_X1 port map( A1 => n147, A2 => n83, ZN => ab_1_29_port);
   U477 : NOR2_X1 port map( A1 => n148, A2 => n83, ZN => ab_1_28_port);
   U478 : NOR2_X1 port map( A1 => n149, A2 => n83, ZN => ab_1_27_port);
   U479 : NOR2_X1 port map( A1 => n150, A2 => n83, ZN => ab_1_26_port);
   U480 : NOR2_X1 port map( A1 => n151, A2 => n83, ZN => ab_1_25_port);
   U481 : NOR2_X1 port map( A1 => n152, A2 => n83, ZN => ab_1_24_port);
   U482 : NOR2_X1 port map( A1 => n153, A2 => n83, ZN => ab_1_23_port);
   U483 : NOR2_X1 port map( A1 => n154, A2 => n83, ZN => ab_1_22_port);
   U484 : NOR2_X1 port map( A1 => n155, A2 => n83, ZN => ab_1_21_port);
   U485 : NOR2_X1 port map( A1 => n156, A2 => n83, ZN => ab_1_20_port);
   U486 : NOR2_X1 port map( A1 => n108, A2 => n82, ZN => ab_1_1_port);
   U487 : NOR2_X1 port map( A1 => n157, A2 => n82, ZN => ab_1_19_port);
   U488 : NOR2_X1 port map( A1 => n158, A2 => n82, ZN => ab_1_18_port);
   U489 : NOR2_X1 port map( A1 => n159, A2 => n82, ZN => ab_1_17_port);
   U490 : NOR2_X1 port map( A1 => n160, A2 => n82, ZN => ab_1_16_port);
   U491 : NOR2_X1 port map( A1 => n161, A2 => n82, ZN => ab_1_15_port);
   U492 : NOR2_X1 port map( A1 => n162, A2 => n82, ZN => ab_1_14_port);
   U493 : NOR2_X1 port map( A1 => n163, A2 => n82, ZN => ab_1_13_port);
   U494 : NOR2_X1 port map( A1 => n164, A2 => n82, ZN => ab_1_12_port);
   U495 : NOR2_X1 port map( A1 => n165, A2 => n82, ZN => ab_1_11_port);
   U496 : NOR2_X1 port map( A1 => n166, A2 => n82, ZN => ab_1_10_port);
   U497 : NOR2_X1 port map( A1 => n111, A2 => n82, ZN => ab_1_0_port);
   U498 : NOR2_X1 port map( A1 => n167, A2 => n125, ZN => ab_19_9_port);
   U499 : NOR2_X1 port map( A1 => n89, A2 => n125, ZN => ab_19_8_port);
   U500 : NOR2_X1 port map( A1 => n91, A2 => n125, ZN => ab_19_7_port);
   U501 : NOR2_X1 port map( A1 => n93, A2 => n125, ZN => ab_19_6_port);
   U502 : NOR2_X1 port map( A1 => n96, A2 => n125, ZN => ab_19_5_port);
   U503 : NOR2_X1 port map( A1 => n99, A2 => n125, ZN => ab_19_4_port);
   U504 : NOR2_X1 port map( A1 => n102, A2 => n125, ZN => ab_19_3_port);
   U505 : NOR2_X1 port map( A1 => n105, A2 => n125, ZN => ab_19_2_port);
   U506 : NOR2_X1 port map( A1 => n108, A2 => n125, ZN => ab_19_1_port);
   U507 : NOR2_X1 port map( A1 => n164, A2 => n125, ZN => ab_19_12_port);
   U508 : NOR2_X1 port map( A1 => n165, A2 => n125, ZN => ab_19_11_port);
   U509 : NOR2_X1 port map( A1 => n166, A2 => n125, ZN => ab_19_10_port);
   U510 : NOR2_X1 port map( A1 => n111, A2 => n125, ZN => ab_19_0_port);
   U511 : NOR2_X1 port map( A1 => n167, A2 => n126, ZN => ab_18_9_port);
   U512 : NOR2_X1 port map( A1 => n89, A2 => n126, ZN => ab_18_8_port);
   U513 : NOR2_X1 port map( A1 => n91, A2 => n126, ZN => ab_18_7_port);
   U514 : NOR2_X1 port map( A1 => n93, A2 => n126, ZN => ab_18_6_port);
   U515 : NOR2_X1 port map( A1 => n96, A2 => n126, ZN => ab_18_5_port);
   U516 : NOR2_X1 port map( A1 => n99, A2 => n126, ZN => ab_18_4_port);
   U517 : NOR2_X1 port map( A1 => n102, A2 => n126, ZN => ab_18_3_port);
   U518 : NOR2_X1 port map( A1 => n105, A2 => n126, ZN => ab_18_2_port);
   U519 : NOR2_X1 port map( A1 => n108, A2 => n126, ZN => ab_18_1_port);
   U520 : NOR2_X1 port map( A1 => n163, A2 => n126, ZN => ab_18_13_port);
   U521 : NOR2_X1 port map( A1 => n164, A2 => n126, ZN => ab_18_12_port);
   U522 : NOR2_X1 port map( A1 => n165, A2 => n126, ZN => ab_18_11_port);
   U523 : NOR2_X1 port map( A1 => n166, A2 => n126, ZN => ab_18_10_port);
   U524 : NOR2_X1 port map( A1 => n111, A2 => n126, ZN => ab_18_0_port);
   U525 : NOR2_X1 port map( A1 => n167, A2 => n127, ZN => ab_17_9_port);
   U526 : NOR2_X1 port map( A1 => n89, A2 => n127, ZN => ab_17_8_port);
   U527 : NOR2_X1 port map( A1 => n91, A2 => n127, ZN => ab_17_7_port);
   U528 : NOR2_X1 port map( A1 => n93, A2 => n127, ZN => ab_17_6_port);
   U529 : NOR2_X1 port map( A1 => n96, A2 => n127, ZN => ab_17_5_port);
   U530 : NOR2_X1 port map( A1 => n99, A2 => n127, ZN => ab_17_4_port);
   U531 : NOR2_X1 port map( A1 => n102, A2 => n127, ZN => ab_17_3_port);
   U532 : NOR2_X1 port map( A1 => n105, A2 => n127, ZN => ab_17_2_port);
   U533 : NOR2_X1 port map( A1 => n108, A2 => n127, ZN => ab_17_1_port);
   U534 : NOR2_X1 port map( A1 => n162, A2 => n127, ZN => ab_17_14_port);
   U535 : NOR2_X1 port map( A1 => n163, A2 => n127, ZN => ab_17_13_port);
   U536 : NOR2_X1 port map( A1 => n164, A2 => n127, ZN => ab_17_12_port);
   U537 : NOR2_X1 port map( A1 => n165, A2 => n127, ZN => ab_17_11_port);
   U538 : NOR2_X1 port map( A1 => n166, A2 => n127, ZN => ab_17_10_port);
   U539 : NOR2_X1 port map( A1 => n111, A2 => n127, ZN => ab_17_0_port);
   U540 : NOR2_X1 port map( A1 => n167, A2 => n128, ZN => ab_16_9_port);
   U541 : NOR2_X1 port map( A1 => n89, A2 => n128, ZN => ab_16_8_port);
   U542 : NOR2_X1 port map( A1 => n91, A2 => n128, ZN => ab_16_7_port);
   U543 : NOR2_X1 port map( A1 => n93, A2 => n128, ZN => ab_16_6_port);
   U544 : NOR2_X1 port map( A1 => n96, A2 => n128, ZN => ab_16_5_port);
   U545 : NOR2_X1 port map( A1 => n99, A2 => n128, ZN => ab_16_4_port);
   U546 : NOR2_X1 port map( A1 => n102, A2 => n128, ZN => ab_16_3_port);
   U547 : NOR2_X1 port map( A1 => n105, A2 => n128, ZN => ab_16_2_port);
   U548 : NOR2_X1 port map( A1 => n108, A2 => n128, ZN => ab_16_1_port);
   U549 : NOR2_X1 port map( A1 => n161, A2 => n128, ZN => ab_16_15_port);
   U550 : NOR2_X1 port map( A1 => n162, A2 => n128, ZN => ab_16_14_port);
   U551 : NOR2_X1 port map( A1 => n163, A2 => n128, ZN => ab_16_13_port);
   U552 : NOR2_X1 port map( A1 => n164, A2 => n128, ZN => ab_16_12_port);
   U553 : NOR2_X1 port map( A1 => n165, A2 => n128, ZN => ab_16_11_port);
   U554 : NOR2_X1 port map( A1 => n166, A2 => n128, ZN => ab_16_10_port);
   U555 : NOR2_X1 port map( A1 => n112, A2 => n128, ZN => ab_16_0_port);
   U556 : NOR2_X1 port map( A1 => n167, A2 => n129, ZN => ab_15_9_port);
   U557 : NOR2_X1 port map( A1 => n89, A2 => n129, ZN => ab_15_8_port);
   U558 : NOR2_X1 port map( A1 => n91, A2 => n129, ZN => ab_15_7_port);
   U559 : NOR2_X1 port map( A1 => n93, A2 => n129, ZN => ab_15_6_port);
   U560 : NOR2_X1 port map( A1 => n96, A2 => n129, ZN => ab_15_5_port);
   U561 : NOR2_X1 port map( A1 => n99, A2 => n129, ZN => ab_15_4_port);
   U562 : NOR2_X1 port map( A1 => n102, A2 => n129, ZN => ab_15_3_port);
   U563 : NOR2_X1 port map( A1 => n105, A2 => n129, ZN => ab_15_2_port);
   U564 : NOR2_X1 port map( A1 => n109, A2 => n129, ZN => ab_15_1_port);
   U565 : NOR2_X1 port map( A1 => n160, A2 => n129, ZN => ab_15_16_port);
   U566 : NOR2_X1 port map( A1 => n161, A2 => n129, ZN => ab_15_15_port);
   U567 : NOR2_X1 port map( A1 => n162, A2 => n129, ZN => ab_15_14_port);
   U568 : NOR2_X1 port map( A1 => n163, A2 => n129, ZN => ab_15_13_port);
   U569 : NOR2_X1 port map( A1 => n164, A2 => n129, ZN => ab_15_12_port);
   U570 : NOR2_X1 port map( A1 => n165, A2 => n129, ZN => ab_15_11_port);
   U571 : NOR2_X1 port map( A1 => n166, A2 => n129, ZN => ab_15_10_port);
   U572 : NOR2_X1 port map( A1 => n112, A2 => n129, ZN => ab_15_0_port);
   U573 : NOR2_X1 port map( A1 => n167, A2 => n130, ZN => ab_14_9_port);
   U574 : NOR2_X1 port map( A1 => n89, A2 => n130, ZN => ab_14_8_port);
   U575 : NOR2_X1 port map( A1 => n91, A2 => n130, ZN => ab_14_7_port);
   U576 : NOR2_X1 port map( A1 => n93, A2 => n130, ZN => ab_14_6_port);
   U577 : NOR2_X1 port map( A1 => n96, A2 => n130, ZN => ab_14_5_port);
   U578 : NOR2_X1 port map( A1 => n99, A2 => n130, ZN => ab_14_4_port);
   U579 : NOR2_X1 port map( A1 => n102, A2 => n130, ZN => ab_14_3_port);
   U580 : NOR2_X1 port map( A1 => n106, A2 => n130, ZN => ab_14_2_port);
   U581 : NOR2_X1 port map( A1 => n109, A2 => n130, ZN => ab_14_1_port);
   U582 : NOR2_X1 port map( A1 => n159, A2 => n130, ZN => ab_14_17_port);
   U583 : NOR2_X1 port map( A1 => n160, A2 => n130, ZN => ab_14_16_port);
   U584 : NOR2_X1 port map( A1 => n161, A2 => n130, ZN => ab_14_15_port);
   U585 : NOR2_X1 port map( A1 => n162, A2 => n130, ZN => ab_14_14_port);
   U586 : NOR2_X1 port map( A1 => n163, A2 => n130, ZN => ab_14_13_port);
   U587 : NOR2_X1 port map( A1 => n164, A2 => n130, ZN => ab_14_12_port);
   U588 : NOR2_X1 port map( A1 => n165, A2 => n130, ZN => ab_14_11_port);
   U589 : NOR2_X1 port map( A1 => n166, A2 => n130, ZN => ab_14_10_port);
   U590 : NOR2_X1 port map( A1 => n112, A2 => n130, ZN => ab_14_0_port);
   U591 : NOR2_X1 port map( A1 => n167, A2 => n131, ZN => ab_13_9_port);
   U592 : NOR2_X1 port map( A1 => n89, A2 => n131, ZN => ab_13_8_port);
   U593 : NOR2_X1 port map( A1 => n91, A2 => n131, ZN => ab_13_7_port);
   U594 : NOR2_X1 port map( A1 => n93, A2 => n131, ZN => ab_13_6_port);
   U595 : NOR2_X1 port map( A1 => n96, A2 => n131, ZN => ab_13_5_port);
   U596 : NOR2_X1 port map( A1 => n99, A2 => n131, ZN => ab_13_4_port);
   U597 : NOR2_X1 port map( A1 => n103, A2 => n131, ZN => ab_13_3_port);
   U598 : NOR2_X1 port map( A1 => n106, A2 => n131, ZN => ab_13_2_port);
   U599 : NOR2_X1 port map( A1 => n109, A2 => n131, ZN => ab_13_1_port);
   U600 : NOR2_X1 port map( A1 => n158, A2 => n131, ZN => ab_13_18_port);
   U601 : NOR2_X1 port map( A1 => n159, A2 => n131, ZN => ab_13_17_port);
   U602 : NOR2_X1 port map( A1 => n160, A2 => n131, ZN => ab_13_16_port);
   U603 : NOR2_X1 port map( A1 => n161, A2 => n131, ZN => ab_13_15_port);
   U604 : NOR2_X1 port map( A1 => n162, A2 => n131, ZN => ab_13_14_port);
   U605 : NOR2_X1 port map( A1 => n163, A2 => n131, ZN => ab_13_13_port);
   U606 : NOR2_X1 port map( A1 => n164, A2 => n131, ZN => ab_13_12_port);
   U607 : NOR2_X1 port map( A1 => n165, A2 => n131, ZN => ab_13_11_port);
   U608 : NOR2_X1 port map( A1 => n166, A2 => n131, ZN => ab_13_10_port);
   U609 : NOR2_X1 port map( A1 => n112, A2 => n131, ZN => ab_13_0_port);
   U610 : NOR2_X1 port map( A1 => n167, A2 => n132, ZN => ab_12_9_port);
   U611 : NOR2_X1 port map( A1 => n89, A2 => n132, ZN => ab_12_8_port);
   U612 : NOR2_X1 port map( A1 => n91, A2 => n132, ZN => ab_12_7_port);
   U613 : NOR2_X1 port map( A1 => n93, A2 => n132, ZN => ab_12_6_port);
   U614 : NOR2_X1 port map( A1 => n96, A2 => n132, ZN => ab_12_5_port);
   U615 : NOR2_X1 port map( A1 => n100, A2 => n132, ZN => ab_12_4_port);
   U616 : NOR2_X1 port map( A1 => n103, A2 => n132, ZN => ab_12_3_port);
   U617 : NOR2_X1 port map( A1 => n106, A2 => n132, ZN => ab_12_2_port);
   U618 : NOR2_X1 port map( A1 => n109, A2 => n132, ZN => ab_12_1_port);
   U619 : NOR2_X1 port map( A1 => n157, A2 => n132, ZN => ab_12_19_port);
   U620 : NOR2_X1 port map( A1 => n158, A2 => n132, ZN => ab_12_18_port);
   U621 : NOR2_X1 port map( A1 => n159, A2 => n132, ZN => ab_12_17_port);
   U622 : NOR2_X1 port map( A1 => n160, A2 => n132, ZN => ab_12_16_port);
   U623 : NOR2_X1 port map( A1 => n161, A2 => n132, ZN => ab_12_15_port);
   U624 : NOR2_X1 port map( A1 => n162, A2 => n132, ZN => ab_12_14_port);
   U625 : NOR2_X1 port map( A1 => n163, A2 => n132, ZN => ab_12_13_port);
   U626 : NOR2_X1 port map( A1 => n164, A2 => n132, ZN => ab_12_12_port);
   U627 : NOR2_X1 port map( A1 => n165, A2 => n132, ZN => ab_12_11_port);
   U628 : NOR2_X1 port map( A1 => n166, A2 => n132, ZN => ab_12_10_port);
   U629 : NOR2_X1 port map( A1 => n112, A2 => n132, ZN => ab_12_0_port);
   U630 : NOR2_X1 port map( A1 => n167, A2 => n133, ZN => ab_11_9_port);
   U631 : NOR2_X1 port map( A1 => n89, A2 => n133, ZN => ab_11_8_port);
   U632 : NOR2_X1 port map( A1 => n91, A2 => n133, ZN => ab_11_7_port);
   U633 : NOR2_X1 port map( A1 => n93, A2 => n133, ZN => ab_11_6_port);
   U634 : NOR2_X1 port map( A1 => n97, A2 => n133, ZN => ab_11_5_port);
   U635 : NOR2_X1 port map( A1 => n100, A2 => n133, ZN => ab_11_4_port);
   U636 : NOR2_X1 port map( A1 => n103, A2 => n133, ZN => ab_11_3_port);
   U637 : NOR2_X1 port map( A1 => n106, A2 => n133, ZN => ab_11_2_port);
   U638 : NOR2_X1 port map( A1 => n156, A2 => n133, ZN => ab_11_20_port);
   U639 : NOR2_X1 port map( A1 => n109, A2 => n133, ZN => ab_11_1_port);
   U640 : NOR2_X1 port map( A1 => n157, A2 => n133, ZN => ab_11_19_port);
   U641 : NOR2_X1 port map( A1 => n158, A2 => n133, ZN => ab_11_18_port);
   U642 : NOR2_X1 port map( A1 => n159, A2 => n133, ZN => ab_11_17_port);
   U643 : NOR2_X1 port map( A1 => n160, A2 => n133, ZN => ab_11_16_port);
   U644 : NOR2_X1 port map( A1 => n161, A2 => n133, ZN => ab_11_15_port);
   U645 : NOR2_X1 port map( A1 => n162, A2 => n133, ZN => ab_11_14_port);
   U646 : NOR2_X1 port map( A1 => n163, A2 => n133, ZN => ab_11_13_port);
   U647 : NOR2_X1 port map( A1 => n164, A2 => n133, ZN => ab_11_12_port);
   U648 : NOR2_X1 port map( A1 => n165, A2 => n133, ZN => ab_11_11_port);
   U649 : NOR2_X1 port map( A1 => n166, A2 => n133, ZN => ab_11_10_port);
   U650 : NOR2_X1 port map( A1 => n112, A2 => n133, ZN => ab_11_0_port);
   U651 : NOR2_X1 port map( A1 => n167, A2 => n134, ZN => ab_10_9_port);
   U652 : NOR2_X1 port map( A1 => n89, A2 => n134, ZN => ab_10_8_port);
   U653 : NOR2_X1 port map( A1 => n91, A2 => n134, ZN => ab_10_7_port);
   U654 : NOR2_X1 port map( A1 => n94, A2 => n134, ZN => ab_10_6_port);
   U655 : NOR2_X1 port map( A1 => n97, A2 => n134, ZN => ab_10_5_port);
   U656 : NOR2_X1 port map( A1 => n100, A2 => n134, ZN => ab_10_4_port);
   U657 : NOR2_X1 port map( A1 => n103, A2 => n134, ZN => ab_10_3_port);
   U658 : NOR2_X1 port map( A1 => n106, A2 => n134, ZN => ab_10_2_port);
   U659 : NOR2_X1 port map( A1 => n155, A2 => n134, ZN => ab_10_21_port);
   U660 : NOR2_X1 port map( A1 => n156, A2 => n134, ZN => ab_10_20_port);
   U661 : NOR2_X1 port map( A1 => n109, A2 => n134, ZN => ab_10_1_port);
   U662 : NOR2_X1 port map( A1 => n157, A2 => n134, ZN => ab_10_19_port);
   U663 : NOR2_X1 port map( A1 => n158, A2 => n134, ZN => ab_10_18_port);
   U664 : NOR2_X1 port map( A1 => n159, A2 => n134, ZN => ab_10_17_port);
   U665 : NOR2_X1 port map( A1 => n160, A2 => n134, ZN => ab_10_16_port);
   U666 : NOR2_X1 port map( A1 => n161, A2 => n134, ZN => ab_10_15_port);
   U667 : NOR2_X1 port map( A1 => n162, A2 => n134, ZN => ab_10_14_port);
   U668 : NOR2_X1 port map( A1 => n163, A2 => n134, ZN => ab_10_13_port);
   U669 : NOR2_X1 port map( A1 => n164, A2 => n134, ZN => ab_10_12_port);
   U670 : NOR2_X1 port map( A1 => n165, A2 => n134, ZN => ab_10_11_port);
   U671 : NOR2_X1 port map( A1 => n166, A2 => n134, ZN => ab_10_10_port);
   U672 : NOR2_X1 port map( A1 => n112, A2 => n134, ZN => ab_10_0_port);
   U673 : NOR2_X1 port map( A1 => n167, A2 => n87, ZN => ab_0_9_port);
   U674 : NOR2_X1 port map( A1 => n89, A2 => n87, ZN => ab_0_8_port);
   U675 : NOR2_X1 port map( A1 => n90, A2 => n87, ZN => ab_0_7_port);
   U676 : NOR2_X1 port map( A1 => n94, A2 => n87, ZN => ab_0_6_port);
   U677 : NOR2_X1 port map( A1 => n97, A2 => n87, ZN => ab_0_5_port);
   U678 : NOR2_X1 port map( A1 => n100, A2 => n87, ZN => ab_0_4_port);
   U679 : NOR2_X1 port map( A1 => n103, A2 => n87, ZN => ab_0_3_port);
   U680 : NOR2_X1 port map( A1 => n145, A2 => n87, ZN => ab_0_31_port);
   U681 : NOR2_X1 port map( A1 => n146, A2 => n86, ZN => ab_0_30_port);
   U682 : NOR2_X1 port map( A1 => n106, A2 => n86, ZN => ab_0_2_port);
   U683 : NOR2_X1 port map( A1 => n147, A2 => n86, ZN => ab_0_29_port);
   U684 : NOR2_X1 port map( A1 => n148, A2 => n86, ZN => ab_0_28_port);
   U685 : NOR2_X1 port map( A1 => n149, A2 => n86, ZN => ab_0_27_port);
   U686 : NOR2_X1 port map( A1 => n150, A2 => n86, ZN => ab_0_26_port);
   U687 : NOR2_X1 port map( A1 => n151, A2 => n86, ZN => ab_0_25_port);
   U688 : NOR2_X1 port map( A1 => n152, A2 => n86, ZN => ab_0_24_port);
   U689 : NOR2_X1 port map( A1 => n153, A2 => n86, ZN => ab_0_23_port);
   U690 : NOR2_X1 port map( A1 => n154, A2 => n86, ZN => ab_0_22_port);
   U691 : NOR2_X1 port map( A1 => n155, A2 => n86, ZN => ab_0_21_port);
   U692 : NOR2_X1 port map( A1 => n156, A2 => n86, ZN => ab_0_20_port);
   U693 : NOR2_X1 port map( A1 => n109, A2 => n85, ZN => ab_0_1_port);
   U694 : NOR2_X1 port map( A1 => n157, A2 => n85, ZN => ab_0_19_port);
   U695 : NOR2_X1 port map( A1 => n158, A2 => n85, ZN => ab_0_18_port);
   U696 : NOR2_X1 port map( A1 => n159, A2 => n85, ZN => ab_0_17_port);
   U697 : NOR2_X1 port map( A1 => n160, A2 => n85, ZN => ab_0_16_port);
   U698 : NOR2_X1 port map( A1 => n161, A2 => n85, ZN => ab_0_15_port);
   U699 : NOR2_X1 port map( A1 => n162, A2 => n85, ZN => ab_0_14_port);
   U700 : NOR2_X1 port map( A1 => n163, A2 => n85, ZN => ab_0_13_port);
   U701 : NOR2_X1 port map( A1 => n164, A2 => n85, ZN => ab_0_12_port);
   U702 : NOR2_X1 port map( A1 => n165, A2 => n85, ZN => ab_0_11_port);
   U703 : NOR2_X1 port map( A1 => n166, A2 => n85, ZN => ab_0_10_port);
   U704 : NOR2_X1 port map( A1 => n112, A2 => n85, ZN => PRODUCT(0));

end SYN_csa;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ALU_ENTITY.all;

entity ALU_ENTITY_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end ALU_ENTITY_DW01_add_0;

architecture SYN_rpl of ALU_ENTITY_DW01_add_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n1, n_1065 : std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1065, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U1 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n1);
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ALU_ENTITY.all;

entity ALU_ENTITY_DW01_sub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end ALU_ENTITY_DW01_sub_0;

architecture SYN_rpl of ALU_ENTITY_DW01_sub_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n1, n2, n3, n4, 
      n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20
      , n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n_1068
      : std_logic;

begin
   
   U2_31 : FA_X1 port map( A => A(31), B => n2, CI => carry_31_port, CO => 
                           n_1068, S => DIFF(31));
   U2_30 : FA_X1 port map( A => A(30), B => n3, CI => carry_30_port, CO => 
                           carry_31_port, S => DIFF(30));
   U2_29 : FA_X1 port map( A => A(29), B => n4, CI => carry_29_port, CO => 
                           carry_30_port, S => DIFF(29));
   U2_28 : FA_X1 port map( A => A(28), B => n5, CI => carry_28_port, CO => 
                           carry_29_port, S => DIFF(28));
   U2_27 : FA_X1 port map( A => A(27), B => n6, CI => carry_27_port, CO => 
                           carry_28_port, S => DIFF(27));
   U2_26 : FA_X1 port map( A => A(26), B => n7, CI => carry_26_port, CO => 
                           carry_27_port, S => DIFF(26));
   U2_25 : FA_X1 port map( A => A(25), B => n8, CI => carry_25_port, CO => 
                           carry_26_port, S => DIFF(25));
   U2_24 : FA_X1 port map( A => A(24), B => n9, CI => carry_24_port, CO => 
                           carry_25_port, S => DIFF(24));
   U2_23 : FA_X1 port map( A => A(23), B => n10, CI => carry_23_port, CO => 
                           carry_24_port, S => DIFF(23));
   U2_22 : FA_X1 port map( A => A(22), B => n11, CI => carry_22_port, CO => 
                           carry_23_port, S => DIFF(22));
   U2_21 : FA_X1 port map( A => A(21), B => n12, CI => carry_21_port, CO => 
                           carry_22_port, S => DIFF(21));
   U2_20 : FA_X1 port map( A => A(20), B => n13, CI => carry_20_port, CO => 
                           carry_21_port, S => DIFF(20));
   U2_19 : FA_X1 port map( A => A(19), B => n14, CI => carry_19_port, CO => 
                           carry_20_port, S => DIFF(19));
   U2_18 : FA_X1 port map( A => A(18), B => n15, CI => carry_18_port, CO => 
                           carry_19_port, S => DIFF(18));
   U2_17 : FA_X1 port map( A => A(17), B => n16, CI => carry_17_port, CO => 
                           carry_18_port, S => DIFF(17));
   U2_16 : FA_X1 port map( A => A(16), B => n17, CI => carry_16_port, CO => 
                           carry_17_port, S => DIFF(16));
   U2_15 : FA_X1 port map( A => A(15), B => n18, CI => carry_15_port, CO => 
                           carry_16_port, S => DIFF(15));
   U2_14 : FA_X1 port map( A => A(14), B => n19, CI => carry_14_port, CO => 
                           carry_15_port, S => DIFF(14));
   U2_13 : FA_X1 port map( A => A(13), B => n20, CI => carry_13_port, CO => 
                           carry_14_port, S => DIFF(13));
   U2_12 : FA_X1 port map( A => A(12), B => n21, CI => carry_12_port, CO => 
                           carry_13_port, S => DIFF(12));
   U2_11 : FA_X1 port map( A => A(11), B => n22, CI => carry_11_port, CO => 
                           carry_12_port, S => DIFF(11));
   U2_10 : FA_X1 port map( A => A(10), B => n23, CI => carry_10_port, CO => 
                           carry_11_port, S => DIFF(10));
   U2_9 : FA_X1 port map( A => A(9), B => n24, CI => carry_9_port, CO => 
                           carry_10_port, S => DIFF(9));
   U2_8 : FA_X1 port map( A => A(8), B => n25, CI => carry_8_port, CO => 
                           carry_9_port, S => DIFF(8));
   U2_7 : FA_X1 port map( A => A(7), B => n26, CI => carry_7_port, CO => 
                           carry_8_port, S => DIFF(7));
   U2_6 : FA_X1 port map( A => A(6), B => n27, CI => carry_6_port, CO => 
                           carry_7_port, S => DIFF(6));
   U2_5 : FA_X1 port map( A => A(5), B => n28, CI => carry_5_port, CO => 
                           carry_6_port, S => DIFF(5));
   U2_4 : FA_X1 port map( A => A(4), B => n29, CI => carry_4_port, CO => 
                           carry_5_port, S => DIFF(4));
   U2_3 : FA_X1 port map( A => A(3), B => n30, CI => carry_3_port, CO => 
                           carry_4_port, S => DIFF(3));
   U2_2 : FA_X1 port map( A => A(2), B => n31, CI => carry_2_port, CO => 
                           carry_3_port, S => DIFF(2));
   U2_1 : FA_X1 port map( A => A(1), B => n32, CI => carry_1_port, CO => 
                           carry_2_port, S => DIFF(1));
   U1 : INV_X1 port map( A => B(31), ZN => n2);
   U2 : INV_X1 port map( A => B(1), ZN => n32);
   U3 : INV_X1 port map( A => A(0), ZN => n1);
   U4 : INV_X1 port map( A => B(2), ZN => n31);
   U5 : INV_X1 port map( A => B(3), ZN => n30);
   U6 : INV_X1 port map( A => B(4), ZN => n29);
   U7 : INV_X1 port map( A => B(5), ZN => n28);
   U8 : INV_X1 port map( A => B(6), ZN => n27);
   U9 : INV_X1 port map( A => B(7), ZN => n26);
   U10 : INV_X1 port map( A => B(8), ZN => n25);
   U11 : INV_X1 port map( A => B(9), ZN => n24);
   U12 : INV_X1 port map( A => B(10), ZN => n23);
   U13 : INV_X1 port map( A => B(11), ZN => n22);
   U14 : INV_X1 port map( A => B(12), ZN => n21);
   U15 : INV_X1 port map( A => B(13), ZN => n20);
   U16 : INV_X1 port map( A => B(14), ZN => n19);
   U17 : INV_X1 port map( A => B(15), ZN => n18);
   U18 : INV_X1 port map( A => B(16), ZN => n17);
   U19 : INV_X1 port map( A => B(17), ZN => n16);
   U20 : INV_X1 port map( A => B(18), ZN => n15);
   U21 : INV_X1 port map( A => B(19), ZN => n14);
   U22 : INV_X1 port map( A => B(20), ZN => n13);
   U23 : INV_X1 port map( A => B(21), ZN => n12);
   U24 : INV_X1 port map( A => B(22), ZN => n11);
   U25 : INV_X1 port map( A => B(23), ZN => n10);
   U26 : INV_X1 port map( A => B(24), ZN => n9);
   U27 : INV_X1 port map( A => B(25), ZN => n8);
   U28 : INV_X1 port map( A => B(26), ZN => n7);
   U29 : INV_X1 port map( A => B(27), ZN => n6);
   U30 : INV_X1 port map( A => B(28), ZN => n5);
   U31 : INV_X1 port map( A => B(29), ZN => n4);
   U32 : INV_X1 port map( A => B(30), ZN => n3);
   U33 : INV_X1 port map( A => B(0), ZN => n33);
   U34 : XNOR2_X1 port map( A => n33, B => A(0), ZN => DIFF(0));
   U35 : NAND2_X1 port map( A1 => B(0), A2 => n1, ZN => carry_1_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ALU_ENTITY.all;

entity ALU_ENTITY is

   port( CLK, RESET : in std_logic;  IN0, IN1 : in std_logic_vector (31 downto 
         0);  OP : in std_logic_vector (2 downto 0);  RESULT : out 
         std_logic_vector (31 downto 0));

end ALU_ENTITY;

architecture SYN_ALU_ARCH of ALU_ENTITY is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component ALU_ENTITY_DW02_mult_0
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  
            PRODUCT : out std_logic_vector (63 downto 0));
   end component;
   
   component ALU_ENTITY_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component ALU_ENTITY_DW01_sub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
      N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58
      , N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, 
      N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87
      , N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
      N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, 
      N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, 
      N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, 
      N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, 
      N278, N279, N280, N281, N282, N283, N284, N285, n1, n2, n40_port, 
      n41_port, n42_port, n43_port, n44_port, n45_port, n46_port, n47_port, 
      n48_port, n49_port, n50_port, n51_port, n52_port, n53_port, n54_port, 
      n55_port, n56_port, n57_port, n58_port, n59_port, n60_port, n61_port, 
      n62_port, n63_port, n64_port, n65_port, n66_port, n67_port, n68_port, 
      n69_port, n70_port, n71_port, n72_port, n73_port, n74_port, n75_port, 
      n76_port, n77_port, n78_port, n79_port, n80_port, n81_port, n82_port, 
      n83_port, n84_port, n85_port, n86_port, n87_port, n88_port, n89_port, 
      n90_port, n91_port, n92_port, n93_port, n94_port, n95_port, n96_port, 
      n97_port, n98_port, n99_port, n100_port, n101_port, n102_port, n103_port,
      n104_port, n105_port, n106_port, n107_port, n108_port, n109_port, 
      n110_port, n111_port, n112_port, n113_port, n114_port, n115_port, 
      n116_port, n117_port, n118_port, n119_port, n120_port, n121_port, 
      n122_port, n123_port, n124_port, n125_port, n126, n127, n128, n129, n130,
      n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, 
      n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
      n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, 
      n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, 
      n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
      n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, 
      n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, 
      n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, 
      n227, n228, n229, n230, n231, n232, n233, n_1069, n_1070, n_1071, n_1072,
      n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, 
      n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, 
      n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, 
      n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, 
      n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, 
      n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, 
      n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134 : 
      std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   RESULT_reg_31_inst : DFF_X1 port map( D => N285, CK => CLK, Q => RESULT(31),
                           QN => n_1069);
   RESULT_reg_30_inst : DFF_X1 port map( D => N284, CK => CLK, Q => RESULT(30),
                           QN => n_1070);
   RESULT_reg_29_inst : DFF_X1 port map( D => N283, CK => CLK, Q => RESULT(29),
                           QN => n_1071);
   RESULT_reg_28_inst : DFF_X1 port map( D => N282, CK => CLK, Q => RESULT(28),
                           QN => n_1072);
   RESULT_reg_27_inst : DFF_X1 port map( D => N281, CK => CLK, Q => RESULT(27),
                           QN => n_1073);
   RESULT_reg_26_inst : DFF_X1 port map( D => N280, CK => CLK, Q => RESULT(26),
                           QN => n_1074);
   RESULT_reg_25_inst : DFF_X1 port map( D => N279, CK => CLK, Q => RESULT(25),
                           QN => n_1075);
   RESULT_reg_24_inst : DFF_X1 port map( D => N278, CK => CLK, Q => RESULT(24),
                           QN => n_1076);
   RESULT_reg_23_inst : DFF_X1 port map( D => N277, CK => CLK, Q => RESULT(23),
                           QN => n_1077);
   RESULT_reg_22_inst : DFF_X1 port map( D => N276, CK => CLK, Q => RESULT(22),
                           QN => n_1078);
   RESULT_reg_21_inst : DFF_X1 port map( D => N275, CK => CLK, Q => RESULT(21),
                           QN => n_1079);
   RESULT_reg_20_inst : DFF_X1 port map( D => N274, CK => CLK, Q => RESULT(20),
                           QN => n_1080);
   RESULT_reg_19_inst : DFF_X1 port map( D => N273, CK => CLK, Q => RESULT(19),
                           QN => n_1081);
   RESULT_reg_18_inst : DFF_X1 port map( D => N272, CK => CLK, Q => RESULT(18),
                           QN => n_1082);
   RESULT_reg_17_inst : DFF_X1 port map( D => N271, CK => CLK, Q => RESULT(17),
                           QN => n_1083);
   RESULT_reg_16_inst : DFF_X1 port map( D => N270, CK => CLK, Q => RESULT(16),
                           QN => n_1084);
   RESULT_reg_15_inst : DFF_X1 port map( D => N269, CK => CLK, Q => RESULT(15),
                           QN => n_1085);
   RESULT_reg_14_inst : DFF_X1 port map( D => N268, CK => CLK, Q => RESULT(14),
                           QN => n_1086);
   RESULT_reg_13_inst : DFF_X1 port map( D => N267, CK => CLK, Q => RESULT(13),
                           QN => n_1087);
   RESULT_reg_12_inst : DFF_X1 port map( D => N266, CK => CLK, Q => RESULT(12),
                           QN => n_1088);
   RESULT_reg_11_inst : DFF_X1 port map( D => N265, CK => CLK, Q => RESULT(11),
                           QN => n_1089);
   RESULT_reg_10_inst : DFF_X1 port map( D => N264, CK => CLK, Q => RESULT(10),
                           QN => n_1090);
   RESULT_reg_9_inst : DFF_X1 port map( D => N263, CK => CLK, Q => RESULT(9), 
                           QN => n_1091);
   RESULT_reg_8_inst : DFF_X1 port map( D => N262, CK => CLK, Q => RESULT(8), 
                           QN => n_1092);
   RESULT_reg_7_inst : DFF_X1 port map( D => N261, CK => CLK, Q => RESULT(7), 
                           QN => n_1093);
   RESULT_reg_6_inst : DFF_X1 port map( D => N260, CK => CLK, Q => RESULT(6), 
                           QN => n_1094);
   RESULT_reg_5_inst : DFF_X1 port map( D => N259, CK => CLK, Q => RESULT(5), 
                           QN => n_1095);
   RESULT_reg_4_inst : DFF_X1 port map( D => N258, CK => CLK, Q => RESULT(4), 
                           QN => n_1096);
   RESULT_reg_3_inst : DFF_X1 port map( D => N257, CK => CLK, Q => RESULT(3), 
                           QN => n_1097);
   RESULT_reg_2_inst : DFF_X1 port map( D => N256, CK => CLK, Q => RESULT(2), 
                           QN => n_1098);
   RESULT_reg_1_inst : DFF_X1 port map( D => N255, CK => CLK, Q => RESULT(1), 
                           QN => n_1099);
   RESULT_reg_0_inst : DFF_X1 port map( D => N254, CK => CLK, Q => RESULT(0), 
                           QN => n_1100);
   U203 : NAND3_X1 port map( A1 => n232, A2 => n231, A3 => OP(2), ZN => 
                           n47_port);
   U204 : NAND2_X1 port map( A1 => OP(2), A2 => n231, ZN => n45_port);
   sub_23 : ALU_ENTITY_DW01_sub_0 port map( A(31) => IN0(31), A(30) => IN0(30),
                           A(29) => IN0(29), A(28) => IN0(28), A(27) => IN0(27)
                           , A(26) => IN0(26), A(25) => IN0(25), A(24) => 
                           IN0(24), A(23) => IN0(23), A(22) => IN0(22), A(21) 
                           => IN0(21), A(20) => IN0(20), A(19) => IN0(19), 
                           A(18) => IN0(18), A(17) => IN0(17), A(16) => IN0(16)
                           , A(15) => IN0(15), A(14) => IN0(14), A(13) => 
                           IN0(13), A(12) => IN0(12), A(11) => IN0(11), A(10) 
                           => IN0(10), A(9) => IN0(9), A(8) => IN0(8), A(7) => 
                           IN0(7), A(6) => IN0(6), A(5) => IN0(5), A(4) => 
                           IN0(4), A(3) => IN0(3), A(2) => IN0(2), A(1) => 
                           IN0(1), A(0) => IN0(0), B(31) => IN1(31), B(30) => 
                           IN1(30), B(29) => IN1(29), B(28) => IN1(28), B(27) 
                           => IN1(27), B(26) => IN1(26), B(25) => IN1(25), 
                           B(24) => IN1(24), B(23) => IN1(23), B(22) => IN1(22)
                           , B(21) => IN1(21), B(20) => IN1(20), B(19) => 
                           IN1(19), B(18) => IN1(18), B(17) => IN1(17), B(16) 
                           => IN1(16), B(15) => IN1(15), B(14) => IN1(14), 
                           B(13) => IN1(13), B(12) => IN1(12), B(11) => IN1(11)
                           , B(10) => IN1(10), B(9) => IN1(9), B(8) => IN1(8), 
                           B(7) => IN1(7), B(6) => IN1(6), B(5) => IN1(5), B(4)
                           => IN1(4), B(3) => IN1(3), B(2) => IN1(2), B(1) => 
                           IN1(1), B(0) => IN1(0), CI => n1, DIFF(31) => N93, 
                           DIFF(30) => N92, DIFF(29) => N91, DIFF(28) => N90, 
                           DIFF(27) => N89, DIFF(26) => N88, DIFF(25) => N87, 
                           DIFF(24) => N86, DIFF(23) => N85, DIFF(22) => N84, 
                           DIFF(21) => N83, DIFF(20) => N82, DIFF(19) => N81, 
                           DIFF(18) => N80, DIFF(17) => N79, DIFF(16) => N78, 
                           DIFF(15) => N77, DIFF(14) => N76, DIFF(13) => N75, 
                           DIFF(12) => N74, DIFF(11) => N73, DIFF(10) => N72, 
                           DIFF(9) => N71, DIFF(8) => N70, DIFF(7) => N69, 
                           DIFF(6) => N68, DIFF(5) => N67, DIFF(4) => N66, 
                           DIFF(3) => N65, DIFF(2) => N64, DIFF(1) => N63, 
                           DIFF(0) => N62, CO => n_1101);
   add_22 : ALU_ENTITY_DW01_add_0 port map( A(31) => IN0(31), A(30) => IN0(30),
                           A(29) => IN0(29), A(28) => IN0(28), A(27) => IN0(27)
                           , A(26) => IN0(26), A(25) => IN0(25), A(24) => 
                           IN0(24), A(23) => IN0(23), A(22) => IN0(22), A(21) 
                           => IN0(21), A(20) => IN0(20), A(19) => IN0(19), 
                           A(18) => IN0(18), A(17) => IN0(17), A(16) => IN0(16)
                           , A(15) => IN0(15), A(14) => IN0(14), A(13) => 
                           IN0(13), A(12) => IN0(12), A(11) => IN0(11), A(10) 
                           => IN0(10), A(9) => IN0(9), A(8) => IN0(8), A(7) => 
                           IN0(7), A(6) => IN0(6), A(5) => IN0(5), A(4) => 
                           IN0(4), A(3) => IN0(3), A(2) => IN0(2), A(1) => 
                           IN0(1), A(0) => IN0(0), B(31) => IN1(31), B(30) => 
                           IN1(30), B(29) => IN1(29), B(28) => IN1(28), B(27) 
                           => IN1(27), B(26) => IN1(26), B(25) => IN1(25), 
                           B(24) => IN1(24), B(23) => IN1(23), B(22) => IN1(22)
                           , B(21) => IN1(21), B(20) => IN1(20), B(19) => 
                           IN1(19), B(18) => IN1(18), B(17) => IN1(17), B(16) 
                           => IN1(16), B(15) => IN1(15), B(14) => IN1(14), 
                           B(13) => IN1(13), B(12) => IN1(12), B(11) => IN1(11)
                           , B(10) => IN1(10), B(9) => IN1(9), B(8) => IN1(8), 
                           B(7) => IN1(7), B(6) => IN1(6), B(5) => IN1(5), B(4)
                           => IN1(4), B(3) => IN1(3), B(2) => IN1(2), B(1) => 
                           IN1(1), B(0) => IN1(0), CI => n2, SUM(31) => N61, 
                           SUM(30) => N60, SUM(29) => N59, SUM(28) => N58, 
                           SUM(27) => N57, SUM(26) => N56, SUM(25) => N55, 
                           SUM(24) => N54, SUM(23) => N53, SUM(22) => N52, 
                           SUM(21) => N51, SUM(20) => N50, SUM(19) => N49, 
                           SUM(18) => N48, SUM(17) => N47, SUM(16) => N46, 
                           SUM(15) => N45, SUM(14) => N44, SUM(13) => N43, 
                           SUM(12) => N42, SUM(11) => N41, SUM(10) => N40, 
                           SUM(9) => N39, SUM(8) => N38, SUM(7) => N37, SUM(6) 
                           => N36, SUM(5) => N35, SUM(4) => N34, SUM(3) => N33,
                           SUM(2) => N32, SUM(1) => N31, SUM(0) => N30, CO => 
                           n_1102);
   mult_25 : ALU_ENTITY_DW02_mult_0 port map( A(31) => IN0(31), A(30) => 
                           IN0(30), A(29) => IN0(29), A(28) => IN0(28), A(27) 
                           => IN0(27), A(26) => IN0(26), A(25) => IN0(25), 
                           A(24) => IN0(24), A(23) => IN0(23), A(22) => IN0(22)
                           , A(21) => IN0(21), A(20) => IN0(20), A(19) => 
                           IN0(19), A(18) => IN0(18), A(17) => IN0(17), A(16) 
                           => IN0(16), A(15) => IN0(15), A(14) => IN0(14), 
                           A(13) => IN0(13), A(12) => IN0(12), A(11) => IN0(11)
                           , A(10) => IN0(10), A(9) => IN0(9), A(8) => IN0(8), 
                           A(7) => IN0(7), A(6) => IN0(6), A(5) => IN0(5), A(4)
                           => IN0(4), A(3) => IN0(3), A(2) => IN0(2), A(1) => 
                           IN0(1), A(0) => IN0(0), B(31) => IN1(31), B(30) => 
                           IN1(30), B(29) => IN1(29), B(28) => IN1(28), B(27) 
                           => IN1(27), B(26) => IN1(26), B(25) => IN1(25), 
                           B(24) => IN1(24), B(23) => IN1(23), B(22) => IN1(22)
                           , B(21) => IN1(21), B(20) => IN1(20), B(19) => 
                           IN1(19), B(18) => IN1(18), B(17) => IN1(17), B(16) 
                           => IN1(16), B(15) => IN1(15), B(14) => IN1(14), 
                           B(13) => IN1(13), B(12) => IN1(12), B(11) => IN1(11)
                           , B(10) => IN1(10), B(9) => IN1(9), B(8) => IN1(8), 
                           B(7) => IN1(7), B(6) => IN1(6), B(5) => IN1(5), B(4)
                           => IN1(4), B(3) => IN1(3), B(2) => IN1(2), B(1) => 
                           IN1(1), B(0) => IN1(0), TC => n233, PRODUCT(63) => 
                           n_1103, PRODUCT(62) => n_1104, PRODUCT(61) => n_1105
                           , PRODUCT(60) => n_1106, PRODUCT(59) => n_1107, 
                           PRODUCT(58) => n_1108, PRODUCT(57) => n_1109, 
                           PRODUCT(56) => n_1110, PRODUCT(55) => n_1111, 
                           PRODUCT(54) => n_1112, PRODUCT(53) => n_1113, 
                           PRODUCT(52) => n_1114, PRODUCT(51) => n_1115, 
                           PRODUCT(50) => n_1116, PRODUCT(49) => n_1117, 
                           PRODUCT(48) => n_1118, PRODUCT(47) => n_1119, 
                           PRODUCT(46) => n_1120, PRODUCT(45) => n_1121, 
                           PRODUCT(44) => n_1122, PRODUCT(43) => n_1123, 
                           PRODUCT(42) => n_1124, PRODUCT(41) => n_1125, 
                           PRODUCT(40) => n_1126, PRODUCT(39) => n_1127, 
                           PRODUCT(38) => n_1128, PRODUCT(37) => n_1129, 
                           PRODUCT(36) => n_1130, PRODUCT(35) => n_1131, 
                           PRODUCT(34) => n_1132, PRODUCT(33) => n_1133, 
                           PRODUCT(32) => n_1134, PRODUCT(31) => N125, 
                           PRODUCT(30) => N124, PRODUCT(29) => N123, 
                           PRODUCT(28) => N122, PRODUCT(27) => N121, 
                           PRODUCT(26) => N120, PRODUCT(25) => N119, 
                           PRODUCT(24) => N118, PRODUCT(23) => N117, 
                           PRODUCT(22) => N116, PRODUCT(21) => N115, 
                           PRODUCT(20) => N114, PRODUCT(19) => N113, 
                           PRODUCT(18) => N112, PRODUCT(17) => N111, 
                           PRODUCT(16) => N110, PRODUCT(15) => N109, 
                           PRODUCT(14) => N108, PRODUCT(13) => N107, 
                           PRODUCT(12) => N106, PRODUCT(11) => N105, 
                           PRODUCT(10) => N104, PRODUCT(9) => N103, PRODUCT(8) 
                           => N102, PRODUCT(7) => N101, PRODUCT(6) => N100, 
                           PRODUCT(5) => N99, PRODUCT(4) => N98, PRODUCT(3) => 
                           N97, PRODUCT(2) => N96, PRODUCT(1) => N95, 
                           PRODUCT(0) => N94);
   U205 : BUF_X1 port map( A => n48_port, Z => n177);
   U206 : BUF_X1 port map( A => n48_port, Z => n178);
   U207 : BUF_X1 port map( A => n49_port, Z => n174);
   U208 : BUF_X1 port map( A => n49_port, Z => n175);
   U209 : BUF_X1 port map( A => n42_port, Z => n194);
   U210 : BUF_X1 port map( A => n42_port, Z => n193);
   U211 : BUF_X1 port map( A => n45_port, Z => n191);
   U212 : BUF_X1 port map( A => n47_port, Z => n181);
   U213 : BUF_X1 port map( A => n46_port, Z => n183);
   U214 : BUF_X1 port map( A => n47_port, Z => n180);
   U215 : BUF_X1 port map( A => n46_port, Z => n184);
   U216 : BUF_X1 port map( A => n45_port, Z => n186);
   U217 : BUF_X1 port map( A => n45_port, Z => n187);
   U218 : BUF_X1 port map( A => n45_port, Z => n190);
   U219 : BUF_X1 port map( A => n45_port, Z => n189);
   U220 : BUF_X1 port map( A => n45_port, Z => n188);
   U221 : BUF_X1 port map( A => n45_port, Z => n192);
   U222 : BUF_X1 port map( A => n48_port, Z => n179);
   U223 : BUF_X1 port map( A => n49_port, Z => n176);
   U224 : BUF_X1 port map( A => n42_port, Z => n195);
   U225 : BUF_X1 port map( A => n47_port, Z => n182);
   U226 : BUF_X1 port map( A => n46_port, Z => n185);
   U227 : AOI21_X1 port map( B1 => n54_port, B2 => n55_port, A => n196, ZN => 
                           N283);
   U228 : AOI22_X1 port map( A1 => N91, A2 => n179, B1 => N59, B2 => n176, ZN 
                           => n54_port);
   U229 : AOI221_X1 port map( B1 => N123, B2 => n193, C1 => IN1(29), C2 => 
                           n56_port, A => n57_port, ZN => n55_port);
   U230 : OAI221_X1 port map( B1 => IN0(29), B2 => n192, C1 => n185, C2 => n201
                           , A => n180, ZN => n56_port);
   U231 : AOI21_X1 port map( B1 => n50_port, B2 => n51_port, A => n196, ZN => 
                           N284);
   U232 : AOI22_X1 port map( A1 => N92, A2 => n179, B1 => N60, B2 => n176, ZN 
                           => n50_port);
   U233 : AOI221_X1 port map( B1 => N124, B2 => n193, C1 => IN1(30), C2 => 
                           n52_port, A => n53_port, ZN => n51_port);
   U234 : OAI221_X1 port map( B1 => IN0(30), B2 => n192, C1 => n185, C2 => n200
                           , A => n180, ZN => n52_port);
   U235 : AOI21_X1 port map( B1 => n40_port, B2 => n41_port, A => n196, ZN => 
                           N285);
   U236 : AOI22_X1 port map( A1 => N93, A2 => n179, B1 => N61, B2 => n176, ZN 
                           => n40_port);
   U237 : AOI221_X1 port map( B1 => N125, B2 => n193, C1 => IN1(31), C2 => 
                           n43_port, A => n44_port, ZN => n41_port);
   U238 : AOI21_X1 port map( B1 => n78_port, B2 => n79_port, A => n196, ZN => 
                           N277);
   U239 : AOI22_X1 port map( A1 => N85, A2 => n178, B1 => N53, B2 => n175, ZN 
                           => n78_port);
   U240 : AOI222_X1 port map( A1 => N117, A2 => n194, B1 => IN0(23), B2 => 
                           n80_port, C1 => IN1(23), C2 => n81_port, ZN => 
                           n79_port);
   U241 : OAI21_X1 port map( B1 => IN1(23), B2 => n189, A => n181, ZN => 
                           n80_port);
   U242 : AOI21_X1 port map( B1 => n66_port, B2 => n67_port, A => n196, ZN => 
                           N280);
   U243 : AOI22_X1 port map( A1 => N88, A2 => n179, B1 => N56, B2 => n176, ZN 
                           => n66_port);
   U244 : AOI222_X1 port map( A1 => N120, A2 => n195, B1 => IN0(26), B2 => 
                           n68_port, C1 => IN1(26), C2 => n69_port, ZN => 
                           n67_port);
   U245 : OAI21_X1 port map( B1 => IN1(26), B2 => n189, A => n182, ZN => 
                           n68_port);
   U246 : AOI21_X1 port map( B1 => n82_port, B2 => n83_port, A => n196, ZN => 
                           N276);
   U247 : AOI22_X1 port map( A1 => N84, A2 => n178, B1 => N52, B2 => n175, ZN 
                           => n82_port);
   U248 : AOI222_X1 port map( A1 => N116, A2 => n194, B1 => IN0(22), B2 => 
                           n84_port, C1 => IN1(22), C2 => n85_port, ZN => 
                           n83_port);
   U249 : OAI21_X1 port map( B1 => IN1(22), B2 => n189, A => n181, ZN => 
                           n84_port);
   U250 : AOI21_X1 port map( B1 => n74_port, B2 => n75_port, A => n196, ZN => 
                           N278);
   U251 : AOI22_X1 port map( A1 => N86, A2 => n179, B1 => N54, B2 => n176, ZN 
                           => n74_port);
   U252 : AOI222_X1 port map( A1 => N118, A2 => n195, B1 => IN0(24), B2 => 
                           n76_port, C1 => IN1(24), C2 => n77_port, ZN => 
                           n75_port);
   U253 : OAI21_X1 port map( B1 => IN1(24), B2 => n189, A => n181, ZN => 
                           n76_port);
   U254 : AOI21_X1 port map( B1 => n86_port, B2 => n87_port, A => n196, ZN => 
                           N275);
   U255 : AOI22_X1 port map( A1 => N83, A2 => n178, B1 => N51, B2 => n175, ZN 
                           => n86_port);
   U256 : AOI221_X1 port map( B1 => N115, B2 => n193, C1 => IN1(21), C2 => 
                           n88_port, A => n89_port, ZN => n87_port);
   U257 : OAI221_X1 port map( B1 => IN0(21), B2 => n192, C1 => n184, C2 => n209
                           , A => n180, ZN => n88_port);
   U258 : AOI21_X1 port map( B1 => n70_port, B2 => n71_port, A => n196, ZN => 
                           N279);
   U259 : AOI22_X1 port map( A1 => N87, A2 => n179, B1 => N55, B2 => n176, ZN 
                           => n70_port);
   U260 : AOI221_X1 port map( B1 => N119, B2 => n193, C1 => IN1(25), C2 => 
                           n72_port, A => n73_port, ZN => n71_port);
   U261 : OAI221_X1 port map( B1 => IN0(25), B2 => n192, C1 => n185, C2 => n205
                           , A => n180, ZN => n72_port);
   U262 : AOI21_X1 port map( B1 => n62_port, B2 => n63_port, A => n196, ZN => 
                           N281);
   U263 : AOI22_X1 port map( A1 => N89, A2 => n179, B1 => N57, B2 => n176, ZN 
                           => n62_port);
   U264 : AOI221_X1 port map( B1 => N121, B2 => n193, C1 => IN1(27), C2 => 
                           n64_port, A => n65_port, ZN => n63_port);
   U265 : OAI221_X1 port map( B1 => IN0(27), B2 => n192, C1 => n185, C2 => n203
                           , A => n180, ZN => n64_port);
   U266 : AOI21_X1 port map( B1 => n58_port, B2 => n59_port, A => n196, ZN => 
                           N282);
   U267 : AOI22_X1 port map( A1 => N90, A2 => n179, B1 => N58, B2 => n176, ZN 
                           => n58_port);
   U268 : AOI221_X1 port map( B1 => N122, B2 => n193, C1 => IN1(28), C2 => 
                           n60_port, A => n61_port, ZN => n59_port);
   U269 : OAI221_X1 port map( B1 => IN0(28), B2 => n192, C1 => n185, C2 => n202
                           , A => n180, ZN => n60_port);
   U270 : AOI21_X1 port map( B1 => n106_port, B2 => n107_port, A => n197, ZN =>
                           N270);
   U271 : AOI22_X1 port map( A1 => N78, A2 => n178, B1 => N46, B2 => n175, ZN 
                           => n106_port);
   U272 : AOI222_X1 port map( A1 => N110, A2 => n194, B1 => IN0(16), B2 => 
                           n108_port, C1 => IN1(16), C2 => n109_port, ZN => 
                           n107_port);
   U273 : OAI21_X1 port map( B1 => IN1(16), B2 => n188, A => n181, ZN => 
                           n108_port);
   U274 : AOI21_X1 port map( B1 => n118_port, B2 => n119_port, A => n197, ZN =>
                           N267);
   U275 : AOI22_X1 port map( A1 => N75, A2 => n178, B1 => N43, B2 => n175, ZN 
                           => n118_port);
   U276 : AOI222_X1 port map( A1 => N107, A2 => n194, B1 => IN0(13), B2 => 
                           n120_port, C1 => IN1(13), C2 => n121_port, ZN => 
                           n119_port);
   U277 : OAI21_X1 port map( B1 => IN1(13), B2 => n188, A => n181, ZN => 
                           n120_port);
   U278 : AOI21_X1 port map( B1 => n114_port, B2 => n115_port, A => n197, ZN =>
                           N268);
   U279 : AOI22_X1 port map( A1 => N76, A2 => n178, B1 => N44, B2 => n175, ZN 
                           => n114_port);
   U280 : AOI222_X1 port map( A1 => N108, A2 => n194, B1 => IN0(14), B2 => 
                           n116_port, C1 => IN1(14), C2 => n117_port, ZN => 
                           n115_port);
   U281 : OAI21_X1 port map( B1 => IN1(14), B2 => n188, A => n181, ZN => 
                           n116_port);
   U282 : AOI21_X1 port map( B1 => n102_port, B2 => n103_port, A => n197, ZN =>
                           N271);
   U283 : AOI22_X1 port map( A1 => N79, A2 => n178, B1 => N47, B2 => n175, ZN 
                           => n102_port);
   U284 : AOI222_X1 port map( A1 => N111, A2 => n194, B1 => IN0(17), B2 => 
                           n104_port, C1 => IN1(17), C2 => n105_port, ZN => 
                           n103_port);
   U285 : OAI21_X1 port map( B1 => IN1(17), B2 => n188, A => n181, ZN => 
                           n104_port);
   U286 : AOI21_X1 port map( B1 => n98_port, B2 => n99_port, A => n197, ZN => 
                           N272);
   U287 : AOI22_X1 port map( A1 => N80, A2 => n178, B1 => N48, B2 => n175, ZN 
                           => n98_port);
   U288 : AOI222_X1 port map( A1 => N112, A2 => n194, B1 => IN0(18), B2 => 
                           n100_port, C1 => IN1(18), C2 => n101_port, ZN => 
                           n99_port);
   U289 : OAI21_X1 port map( B1 => IN1(18), B2 => n189, A => n181, ZN => 
                           n100_port);
   U290 : AOI21_X1 port map( B1 => n110_port, B2 => n111_port, A => n197, ZN =>
                           N269);
   U291 : AOI22_X1 port map( A1 => N77, A2 => n178, B1 => N45, B2 => n175, ZN 
                           => n110_port);
   U292 : AOI221_X1 port map( B1 => N109, B2 => n193, C1 => IN1(15), C2 => 
                           n112_port, A => n113_port, ZN => n111_port);
   U293 : OAI221_X1 port map( B1 => IN0(15), B2 => n191, C1 => n184, C2 => n215
                           , A => n180, ZN => n112_port);
   U294 : AOI21_X1 port map( B1 => n94_port, B2 => n95_port, A => n197, ZN => 
                           N273);
   U295 : AOI22_X1 port map( A1 => N81, A2 => n178, B1 => N49, B2 => n175, ZN 
                           => n94_port);
   U296 : AOI221_X1 port map( B1 => N113, B2 => n193, C1 => IN1(19), C2 => 
                           n96_port, A => n97_port, ZN => n95_port);
   U297 : OAI221_X1 port map( B1 => IN0(19), B2 => n191, C1 => n184, C2 => n211
                           , A => n180, ZN => n96_port);
   U298 : AOI21_X1 port map( B1 => n90_port, B2 => n91_port, A => n196, ZN => 
                           N274);
   U299 : AOI22_X1 port map( A1 => N82, A2 => n178, B1 => N50, B2 => n175, ZN 
                           => n90_port);
   U300 : AOI221_X1 port map( B1 => N114, B2 => n193, C1 => IN1(20), C2 => 
                           n92_port, A => n93_port, ZN => n91_port);
   U301 : OAI221_X1 port map( B1 => IN0(20), B2 => n192, C1 => n184, C2 => n210
                           , A => n180, ZN => n92_port);
   U302 : AOI21_X1 port map( B1 => n150, B2 => n151, A => n198, ZN => N259);
   U303 : AOI22_X1 port map( A1 => N67, A2 => n177, B1 => N35, B2 => n174, ZN 
                           => n150);
   U304 : AOI222_X1 port map( A1 => N99, A2 => n195, B1 => IN0(5), B2 => n152, 
                           C1 => IN1(5), C2 => n153, ZN => n151);
   U305 : OAI21_X1 port map( B1 => IN1(5), B2 => n187, A => n182, ZN => n152);
   U306 : AOI21_X1 port map( B1 => n146, B2 => n147, A => n198, ZN => N260);
   U307 : AOI22_X1 port map( A1 => N68, A2 => n177, B1 => N36, B2 => n174, ZN 
                           => n146);
   U308 : AOI222_X1 port map( A1 => N100, A2 => n195, B1 => IN0(6), B2 => n148,
                           C1 => IN1(6), C2 => n149, ZN => n147);
   U309 : OAI21_X1 port map( B1 => IN1(6), B2 => n187, A => n182, ZN => n148);
   U310 : AOI21_X1 port map( B1 => n142, B2 => n143, A => n198, ZN => N261);
   U311 : AOI22_X1 port map( A1 => N69, A2 => n177, B1 => N37, B2 => n174, ZN 
                           => n142);
   U312 : AOI221_X1 port map( B1 => N101, B2 => n194, C1 => IN1(7), C2 => n144,
                           A => n145, ZN => n143);
   U313 : NOR3_X1 port map( A1 => n223, A2 => IN1(7), A3 => n187, ZN => n145);
   U314 : AOI21_X1 port map( B1 => n134, B2 => n135, A => n197, ZN => N263);
   U315 : AOI22_X1 port map( A1 => N71, A2 => n177, B1 => N39, B2 => n174, ZN 
                           => n134);
   U316 : AOI222_X1 port map( A1 => N103, A2 => n194, B1 => IN0(9), B2 => n136,
                           C1 => IN1(9), C2 => n137, ZN => n135);
   U317 : OAI21_X1 port map( B1 => IN1(9), B2 => n187, A => n181, ZN => n136);
   U318 : AOI21_X1 port map( B1 => n130, B2 => n131, A => n197, ZN => N264);
   U319 : AOI22_X1 port map( A1 => N72, A2 => n177, B1 => N40, B2 => n174, ZN 
                           => n130);
   U320 : AOI222_X1 port map( A1 => N104, A2 => n194, B1 => IN0(10), B2 => n132
                           , C1 => IN1(10), C2 => n133, ZN => n131);
   U321 : OAI21_X1 port map( B1 => IN1(10), B2 => n188, A => n181, ZN => n132);
   U322 : AOI21_X1 port map( B1 => n122_port, B2 => n123_port, A => n197, ZN =>
                           N266);
   U323 : AOI22_X1 port map( A1 => N74, A2 => n178, B1 => N42, B2 => n175, ZN 
                           => n122_port);
   U324 : AOI222_X1 port map( A1 => N106, A2 => n194, B1 => IN0(12), B2 => 
                           n124_port, C1 => IN1(12), C2 => n125_port, ZN => 
                           n123_port);
   U325 : OAI21_X1 port map( B1 => IN1(12), B2 => n188, A => n181, ZN => 
                           n124_port);
   U326 : AOI21_X1 port map( B1 => n138, B2 => n139, A => n197, ZN => N262);
   U327 : AOI22_X1 port map( A1 => N70, A2 => n177, B1 => N38, B2 => n174, ZN 
                           => n138);
   U328 : AOI221_X1 port map( B1 => N102, B2 => n194, C1 => IN1(8), C2 => n140,
                           A => n141, ZN => n139);
   U329 : NOR3_X1 port map( A1 => n222, A2 => IN1(8), A3 => n187, ZN => n141);
   U330 : AOI21_X1 port map( B1 => n126, B2 => n127, A => n197, ZN => N265);
   U331 : AOI22_X1 port map( A1 => N73, A2 => n177, B1 => N41, B2 => n174, ZN 
                           => n126);
   U332 : AOI221_X1 port map( B1 => N105, B2 => n193, C1 => IN1(11), C2 => n128
                           , A => n129, ZN => n127);
   U333 : OAI221_X1 port map( B1 => IN0(11), B2 => n191, C1 => n184, C2 => n219
                           , A => n180, ZN => n128);
   U334 : OAI221_X1 port map( B1 => IN0(7), B2 => n191, C1 => n184, C2 => n223,
                           A => n181, ZN => n144);
   U335 : OAI221_X1 port map( B1 => IN0(8), B2 => n191, C1 => n184, C2 => n222,
                           A => n181, ZN => n140);
   U336 : OAI221_X1 port map( B1 => IN0(0), B2 => n192, C1 => n185, C2 => n230,
                           A => n180, ZN => n172);
   U337 : OAI221_X1 port map( B1 => IN0(31), B2 => n192, C1 => n199, C2 => n183
                           , A => n180, ZN => n43_port);
   U338 : NOR3_X1 port map( A1 => OP(0), A2 => OP(2), A3 => n231, ZN => 
                           n42_port);
   U339 : NOR3_X1 port map( A1 => OP(1), A2 => OP(2), A3 => n232, ZN => 
                           n48_port);
   U340 : NOR3_X1 port map( A1 => OP(1), A2 => OP(2), A3 => OP(0), ZN => 
                           n49_port);
   U341 : OAI22_X1 port map( A1 => n183, A2 => n229, B1 => IN0(1), B2 => n191, 
                           ZN => n169);
   U342 : INV_X1 port map( A => IN0(1), ZN => n229);
   U343 : OAI22_X1 port map( A1 => n183, A2 => n228, B1 => IN0(2), B2 => n191, 
                           ZN => n165);
   U344 : INV_X1 port map( A => IN0(2), ZN => n228);
   U345 : OAI22_X1 port map( A1 => n183, A2 => n214, B1 => IN0(16), B2 => n191,
                           ZN => n109_port);
   U346 : INV_X1 port map( A => IN0(16), ZN => n214);
   U347 : OAI22_X1 port map( A1 => n184, A2 => n207, B1 => IN0(23), B2 => n191,
                           ZN => n81_port);
   U348 : INV_X1 port map( A => IN0(23), ZN => n207);
   U349 : OAI22_X1 port map( A1 => n184, A2 => n204, B1 => IN0(26), B2 => n191,
                           ZN => n69_port);
   U350 : INV_X1 port map( A => IN0(26), ZN => n204);
   U351 : BUF_X1 port map( A => RESET, Z => n197);
   U352 : BUF_X1 port map( A => RESET, Z => n196);
   U353 : OAI22_X1 port map( A1 => n183, A2 => n225, B1 => IN0(5), B2 => n189, 
                           ZN => n153);
   U354 : INV_X1 port map( A => IN0(5), ZN => n225);
   U355 : OAI22_X1 port map( A1 => n183, A2 => n220, B1 => IN0(10), B2 => n189,
                           ZN => n133);
   U356 : INV_X1 port map( A => IN0(10), ZN => n220);
   U357 : OAI22_X1 port map( A1 => n183, A2 => n218, B1 => IN0(12), B2 => n189,
                           ZN => n125_port);
   U358 : INV_X1 port map( A => IN0(12), ZN => n218);
   U359 : OAI22_X1 port map( A1 => n183, A2 => n216, B1 => IN0(14), B2 => n189,
                           ZN => n117_port);
   U360 : INV_X1 port map( A => IN0(14), ZN => n216);
   U361 : OAI22_X1 port map( A1 => n183, A2 => n227, B1 => IN0(3), B2 => n190, 
                           ZN => n161);
   U362 : INV_X1 port map( A => IN0(3), ZN => n227);
   U363 : OAI22_X1 port map( A1 => n183, A2 => n226, B1 => IN0(4), B2 => n190, 
                           ZN => n157);
   U364 : INV_X1 port map( A => IN0(4), ZN => n226);
   U365 : OAI22_X1 port map( A1 => n183, A2 => n224, B1 => IN0(6), B2 => n190, 
                           ZN => n149);
   U366 : INV_X1 port map( A => IN0(6), ZN => n224);
   U367 : OAI22_X1 port map( A1 => n183, A2 => n221, B1 => IN0(9), B2 => n190, 
                           ZN => n137);
   U368 : INV_X1 port map( A => IN0(9), ZN => n221);
   U369 : OAI22_X1 port map( A1 => n183, A2 => n217, B1 => IN0(13), B2 => n190,
                           ZN => n121_port);
   U370 : INV_X1 port map( A => IN0(13), ZN => n217);
   U371 : OAI22_X1 port map( A1 => n184, A2 => n213, B1 => IN0(17), B2 => n190,
                           ZN => n105_port);
   U372 : INV_X1 port map( A => IN0(17), ZN => n213);
   U373 : OAI22_X1 port map( A1 => n184, A2 => n212, B1 => IN0(18), B2 => n190,
                           ZN => n101_port);
   U374 : INV_X1 port map( A => IN0(18), ZN => n212);
   U375 : OAI22_X1 port map( A1 => n184, A2 => n208, B1 => IN0(22), B2 => n190,
                           ZN => n85_port);
   U376 : INV_X1 port map( A => IN0(22), ZN => n208);
   U377 : OAI22_X1 port map( A1 => n184, A2 => n206, B1 => IN0(24), B2 => n190,
                           ZN => n77_port);
   U378 : INV_X1 port map( A => IN0(24), ZN => n206);
   U379 : NOR3_X1 port map( A1 => n230, A2 => IN1(0), A3 => n187, ZN => n173);
   U380 : NOR3_X1 port map( A1 => n219, A2 => IN1(11), A3 => n187, ZN => n129);
   U381 : NOR3_X1 port map( A1 => n215, A2 => IN1(15), A3 => n187, ZN => 
                           n113_port);
   U382 : NOR3_X1 port map( A1 => n211, A2 => IN1(19), A3 => n186, ZN => 
                           n97_port);
   U383 : NOR3_X1 port map( A1 => n210, A2 => IN1(20), A3 => n186, ZN => 
                           n93_port);
   U384 : NOR3_X1 port map( A1 => n209, A2 => IN1(21), A3 => n186, ZN => 
                           n89_port);
   U385 : NOR3_X1 port map( A1 => n205, A2 => IN1(25), A3 => n186, ZN => 
                           n73_port);
   U386 : NOR3_X1 port map( A1 => n203, A2 => IN1(27), A3 => n186, ZN => 
                           n65_port);
   U387 : NOR3_X1 port map( A1 => n202, A2 => IN1(28), A3 => n186, ZN => 
                           n61_port);
   U388 : NOR3_X1 port map( A1 => n201, A2 => IN1(29), A3 => n186, ZN => 
                           n57_port);
   U389 : NOR3_X1 port map( A1 => n200, A2 => IN1(30), A3 => n186, ZN => 
                           n53_port);
   U390 : NOR3_X1 port map( A1 => n199, A2 => IN1(31), A3 => n186, ZN => 
                           n44_port);
   U391 : BUF_X1 port map( A => RESET, Z => n198);
   U392 : INV_X1 port map( A => OP(1), ZN => n231);
   U393 : AOI21_X1 port map( B1 => n170, B2 => n171, A => n198, ZN => N254);
   U394 : AOI22_X1 port map( A1 => N62, A2 => n177, B1 => N30, B2 => n174, ZN 
                           => n170);
   U395 : AOI221_X1 port map( B1 => N94, B2 => n193, C1 => IN1(0), C2 => n172, 
                           A => n173, ZN => n171);
   U396 : AOI21_X1 port map( B1 => n166, B2 => n167, A => n198, ZN => N255);
   U397 : AOI22_X1 port map( A1 => N63, A2 => n177, B1 => N31, B2 => n174, ZN 
                           => n166);
   U398 : AOI222_X1 port map( A1 => N95, A2 => n195, B1 => IN0(1), B2 => n168, 
                           C1 => IN1(1), C2 => n169, ZN => n167);
   U399 : OAI21_X1 port map( B1 => IN1(1), B2 => n188, A => n182, ZN => n168);
   U400 : AOI21_X1 port map( B1 => n162, B2 => n163, A => n198, ZN => N256);
   U401 : AOI22_X1 port map( A1 => N64, A2 => n177, B1 => N32, B2 => n174, ZN 
                           => n162);
   U402 : AOI222_X1 port map( A1 => N96, A2 => n195, B1 => IN0(2), B2 => n164, 
                           C1 => IN1(2), C2 => n165, ZN => n163);
   U403 : OAI21_X1 port map( B1 => IN1(2), B2 => n188, A => n182, ZN => n164);
   U404 : AOI21_X1 port map( B1 => n158, B2 => n159, A => n198, ZN => N257);
   U405 : AOI22_X1 port map( A1 => N65, A2 => n177, B1 => N33, B2 => n174, ZN 
                           => n158);
   U406 : AOI222_X1 port map( A1 => N97, A2 => n195, B1 => IN0(3), B2 => n160, 
                           C1 => IN1(3), C2 => n161, ZN => n159);
   U407 : OAI21_X1 port map( B1 => IN1(3), B2 => n187, A => n182, ZN => n160);
   U408 : AOI21_X1 port map( B1 => n154, B2 => n155, A => n198, ZN => N258);
   U409 : AOI22_X1 port map( A1 => N66, A2 => n177, B1 => N34, B2 => n174, ZN 
                           => n154);
   U410 : AOI222_X1 port map( A1 => N98, A2 => n195, B1 => IN0(4), B2 => n156, 
                           C1 => IN1(4), C2 => n157, ZN => n155);
   U411 : OAI21_X1 port map( B1 => IN1(4), B2 => n188, A => n182, ZN => n156);
   U412 : INV_X1 port map( A => OP(0), ZN => n232);
   U413 : OR3_X1 port map( A1 => n232, A2 => OP(2), A3 => n231, ZN => n46_port)
                           ;
   U414 : INV_X1 port map( A => IN0(0), ZN => n230);
   U415 : INV_X1 port map( A => IN0(7), ZN => n223);
   U416 : INV_X1 port map( A => IN0(8), ZN => n222);
   U417 : INV_X1 port map( A => IN0(11), ZN => n219);
   U418 : INV_X1 port map( A => IN0(15), ZN => n215);
   U419 : INV_X1 port map( A => IN0(19), ZN => n211);
   U420 : INV_X1 port map( A => IN0(20), ZN => n210);
   U421 : INV_X1 port map( A => IN0(21), ZN => n209);
   U422 : INV_X1 port map( A => IN0(25), ZN => n205);
   U423 : INV_X1 port map( A => IN0(27), ZN => n203);
   U424 : INV_X1 port map( A => IN0(28), ZN => n202);
   U425 : INV_X1 port map( A => IN0(29), ZN => n201);
   U426 : INV_X1 port map( A => IN0(30), ZN => n200);
   U427 : INV_X1 port map( A => IN0(31), ZN => n199);
   n233 <= '0';

end SYN_ALU_ARCH;
