LIBRARY IEEE;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.std_logic_1164.ALL;

ENTITY ALU_ENTITY IS
	PORT(CLK, RESET : IN STD_LOGIC;
		IN0,IN1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		OP: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		RESULT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END ENTITY;

ARCHITECTURE ALU_ARCH OF ALU_ENTITY IS
BEGIN
    PROCESS(CLK) 
    VARIABLE TMP : STD_LOGIC_VECTOR(63 DOWNTO 0);
    BEGIN
		IF RISING_EDGE(CLK) THEN
			IF RESET = '1' THEN
				 RESULT <= (OTHERS => '0');
			ELSE
				 CASE(OP) IS
					WHEN "000" => RESULT <= UNSIGNED(IN0) + UNSIGNED(IN1);
					WHEN "001" => RESULT <= UNSIGNED(IN0) - UNSIGNED(IN1);
					WHEN "010" => 
						TMP := UNSIGNED(IN0) * UNSIGNED(IN1);
						RESULT <= TMP(31 DOWNTO 0);
					WHEN "011" => RESULT <= IN0 AND IN1;
					WHEN "100" => RESULT <= IN0 OR IN1;
					WHEN "101" => RESULT <= IN0 XOR IN1;
					WHEN OTHERS => RESULT <= (OTHERS => '0');
				 END CASE;
			END IF;
		END IF;
	END PROCESS;
END ARCHITECTURE;
